///////////////////////////////////////////////////////
//	File Name: adc045_wrap.routed.v
//	Data:      25/04/09 13:22:04
//	Program:   xcore
///////////////////////////////////////////////////////
//
module adc045_wrap ( cs, dout, drdy, hard_start, hard_wreg, rst_l, rst_l_adc, din, nRST, ready_sample, sclk, start, clk,  adc045_data );
  input cs, dout, drdy, hard_start, hard_wreg, rst_l, rst_l_adc, clk;
  output din, nRST, ready_sample, sclk, start;
  output  [23:0] adc045_data;
  wire \net21156<0> , \net8287<5> , \net8296<11> , \net8296<10> , \net8296<5> , \net8299<13> , \net8311<10> , \LongBus_20<5> , \LongBus_20<7> , \net8311<8> , 
    \LongBus_20<2> , \net8311<13> , \LongBus_21<12> , \net8320<3> , \net8320<6> , \LongBus_21<9> , \LongBus_21<11> , \net8320<4> , \net8320<5> , \LongBus_21<10> , 
    \LongBus_21<13> , \net8320<2> , \net8320<7> , \LongBus_21<15> , \net8320<0> , \net8320<1> , \LongBus_21<14> , \LongBus_21<3> , \net8320<12> , \net8320<13> , 
    \LongBus_19<10> , \LongBus_3<11> , \LongBus_3<5> , \LongBus_3<4> , \LongBus_3<1> , \LongBus_2<9> , \LongBus_2<10> , \LongBus_2<4> , \LongBus_2<0> , \LongBus_2<2> , 
    \LongBus_2<3> , \LongBus_2<15> , \LongBus_5<14> , \LongBus_0<14> , \LongBus_0<5> , \LongBus_0<0> , \LongBus_0<1> , \LongBus_0<2> , \LongBus_6<10> , \LongBus_6<5> , 
    \LongBus_6<4> , \LongBus_6<2> , \LongBus_1<8> , \LongBus_1<10> , \LongBus_1<7> , \LongBus_1<5> , \LongBus_1<4> , \LongBus_1<0> , \LongBus_1<1> , \LongBus_1<2> , 
    \I3621.I152.net117 , \net10329<2> , \net9202<2> , \LongBus_68<4> , \LongBus_68<5> , \LongBus_68<2> , \LongBus_69<14> , \LongBus_69<15> , \LongBus_68<3> , \LongBus_79<5> , 
    \LongBus_78<4> , \LongBus_78<5> , \LongBus_78<6> , \LongBus_78<9> , \LongBus_78<10> , \LongBus_78<13> , \LongBus_78<14> , \LongBus_78<3> , \LongBus_78<2> , \LongBus_78<1> , 
    \LongBus_78<0> , \LongBus_73<4> , \LongBus_73<5> , \LongBus_73<12> , \LongBus_73<9> , \LongBus_73<11> , \LongBus_73<10> , \LongBus_73<13> , \LongBus_73<8> , \LongBus_73<15> , 
    \LongBus_73<14> , \LongBus_73<1> , \LongBus_73<0> , \LongBus_72<11> , \LongBus_72<10> , \LongBus_72<14> , \LongBus_72<2> , \LongBus_72<1> , \LongBus_70<4> , \LongBus_70<5> , 
    \LongBus_70<7> , \LongBus_70<2> , \LongBus_70<1> , \LongBus_70<0> , \LongBus_71<4> , \LongBus_71<5> , \LongBus_71<11> , \LongBus_71<15> , \LongBus_71<14> , \LongBus_71<3> , 
    \LongBus_71<2> , \I3590.net66 , \I3590.net052 , \I3590.net72 , \I3590.net059 , \I3590.net78 , \I3590.net84 , \I3590.net073 , \net10305<0> , \net10281<1> , 
    \net10281<0> , \net10305<1> , \net10262<3> , \net10262<2> , \net10262<1> , \net10262<0> , \I3690.net35 , \net20974<3> , \I3690.net39 , \net20974<2> , 
    \I3690.net43 , \net20974<1> , \I3690.net47 , \net20974<0> , \I3689.net35 , \net20977<3> , \I3689.net39 , \net20977<2> , \I3687.net43 , \net21016<1> , 
    \GCLK_s1<0> , \GCLK_s1<1> , \GCLK_s1<2> , \net20955<0> , \net16222<3> , \net16222<2> , \GCLK_s5<2> , \ILAB0102.I5605.net25 , \ILAB0102.Clk_int<1> , \ILAB0102.I5605.net29 , 
    \ILAB0102.Clk_int<3> , \ILAB0102.net027166 , \ILAB0102.net27188 , \ILAB0102.I5366.net64 , \ILAB0102.I5366.net68 , \ILAB0102.I5366.net0114 , \ILAB0102.net15299<3> , \ILAB0102.I5366.net0110 , \ILAB0102.net15299<2> , \ILAB0102.I5366.net0106 , 
    \ILAB0102.net15299<1> , \ILAB0102.I5366.net0102 , \ILAB0102.net15299<0> , \ILAB0102.Clk_LAB<0> , \ILAB0102.Clk_LAB<1> , \ILAB0102.Clk_LAB<2> , \ILAB0102.Clk_LAB<3> , \ILAB0102.net18266 , \ILAB0102.net24386 , \ILAB0102.net15476 , 
    \ILAB0102.net26501 , \ILAB0102.net22001 , \net17151<0> , \ILAB0102.net38382 , \net10350<1> , \ILAB0102.net27291 , \ILAB0102.net38760 , \net10355<1> , \ILAB0102.net27305 , \net17150<0> , 
    \ILAB0102.net39618 , \net17154<0> , \ILAB0102.net38964 , \net10357<1> , \ILAB0102.net27339 , \ILAB0102.net22856 , \ILAB0102.net37425 , \net17149<0> , \ILAB0102.net39222 , \net17152<0> , 
    \ILAB0102.net39858 , \ILAB0102.net39579 , \ILAB0102.net16421 , \ILAB0102.net40197 , \ILAB0102.net26726 , \ILAB0102.net40017 , \ILAB0102.net38148 , \ILAB0102.ILE1607.net0562 , \ILAB0102.net15863 , \net18568<0> , 
    \ILAB0102.net19624 , \Fast_out_28<0> , \ILAB0102.net17527 , \ILAB0102.net25852 , \ILAB0102.net23332 , \ILAB0102.net15367 , \ILAB0102.net16132 , \ILAB0102.net21064 , \ILAB0102.ILE0308.net2656 , \ILAB0102.net18562 , 
    \net18584<1> , \net18584<2> , \ILAB0102.net26482 , \ILAB0102.net15482 , \ILAB0102.net26014 , \ILAB0102.net20182 , \ILAB0102.net20722 , \ILAB0102.net15548 , \ILAB0102.net25609 , \net10426<6> , 
    \Fast_out_28<4> , \ILAB0102.net25020 , \ILAB0102.ILE0404.net2656 , \ILAB0102.net20029 , \ILAB0102.net16652 , \ILAB0102.net16654 , \ILAB0102.net15637 , \ILAB0102.net15817 , \ILAB0102.net17419 , \ILAB0102.net26456 , 
    \net17210<3> , \ILAB0102.net16924 , \ILAB0102.net15709 , \ILAB0102.net20344 , \ILAB0102.net20340 , \ILAB0102.ILE0703.net2656 , \ILAB0102.ILE0703.net0541 , \ILAB0102.net17707 , \ILAB0102.net16177 , \ILAB0102.net26347 , 
    \ILAB0102.net15728 , \ILAB0102.net20857 , \net18576<3> , \ILAB0102.net15754 , \ILAB0102.net15889 , \ILAB0102.ILE1505.net2656 , \ILAB0102.net17374 , \ILAB0102.net25989 , \ILAB0102.net25988 , \ILAB0102.net26392 , 
    \ILAB0102.net17663 , \ILAB0102.net15799 , \ILAB0102.net15844 , \ILAB0102.ILE0605.net2656 , \ILAB0102.net15818 , \ILAB0102.net17959 , \ILAB0102.ILE0705.net2656 , \ILAB0102.ILE1605.net0562 , \ILAB0102.net15864 , \ILAB0102.ILE1605.net2656 , 
    \ILAB0102.net25067 , \ILAB0102.net16627 , \ILAB0102.net25133 , \ILAB0102.net15908 , \ILAB0102.net16628 , \ILAB0102.net15907 , \ILAB0102.net20452 , \ILAB0102.net15934 , \ILAB0102.net25069 , \ILAB0102.net25065 , 
    \ILAB0102.ILE1305.net2656 , \ILAB0102.net18229 , \ILAB0102.net24664 , \ILAB0102.net16069 , \ILAB0102.net18634 , \ILAB0102.ILE0706.net2656 , \ILAB0102.net25114 , \ILAB0102.net26797 , \net17226<6> , \ILAB0102.ILE0304.net2656 , 
    \ILAB0102.net26366 , \ILAB0102.ILE1504.net2656 , \ILAB0102.net17122 , \ILAB0102.net16222 , \ILAB0102.net17032 , \ILAB0102.net16267 , \ILAB0102.net25807 , \ILAB0102.net18202 , \ILAB0102.net17167 , \ILAB0102.net16357 , 
    \ILAB0102.net17932 , \ILAB0102.net19129 , \ILAB0102.net16852 , \ILAB0102.net18407 , \ILAB0102.ILE0309.net2656 , \net17198<6> , \ILAB0102.ILE1001.net01345 , \net17198<1> , \ILAB0102.net16537 , \ILAB0102.net16601 , 
    \net17194<3> , \net17194<6> , \ILAB0102.ILE1101.net01339 , \ILAB0102.ILE1303.net0560 , \ILAB0102.ILE1303.net2656 , \ILAB0102.net18112 , \ILAB0102.net17753 , \ILAB0102.net16672 , \ILAB0102.net25249 , \ILAB0102.net17102 , 
    \ILAB0102.ILE0407.net2656 , \ILAB0102.net25447 , \ILAB0102.net18744 , \ILAB0102.net24997 , \ILAB0102.net16763 , \ILAB0102.net25448 , \ILAB0102.net16762 , \ILAB0102.net25969 , \ILAB0102.ILE0507.net2656 , \ILAB0102.net23827 , 
    \ILAB0102.net26662 , \ILAB0102.ILE1103.net2656 , \net17155<1> , \net17230<6> , \ILAB0102.net20614 , \ILAB0102.net19796 , \ILAB0102.net19309 , \net10423<3> , \ILAB0102.ILE0516.net01339 , \net10423<0> , 
    \net10423<6> , \ILAB0102.net17509 , \ILAB0102.net17014 , \ILAB0102.ILE0516.net2656 , \ILAB0102.net25744 , \ILAB0102.net17149 , \ILAB0102.ILE0607.net2656 , \ILAB0102.net18699 , \ILAB0102.ILE1307.net2656 , \ILAB0102.net17194 , 
    \ILAB0102.net17214 , \ILAB0102.ILE0707.net2656 , \Fast_out_28<2> , \net10358<0> , \net10427<1> , \net10427<3> , \ILAB0102.ILE0416.net0562 , \ILAB0102.ILE0416.net0558 , \net10427<5> , \ILAB0102.net19238 , 
    \ILAB0102.ILE0416.net2656 , \ILAB0102.net25584 , \ILAB0102.net17347 , \ILAB0102.ILE0805.net2656 , \ILAB0102.net26617 , \ILAB0102.ILE1003.net0562 , \ILAB0102.ILE1003.net2656 , \ILAB0102.net21739 , \net10411<1> , \ILAB0102.net18878 , 
    \ILAB0102.net18652 , \ILAB0102.ILE0816.net2656 , \net10407<1> , \ILAB0102.net22164 , \net10407<2> , \net10407<0> , \net10407<6> , \ILAB0102.net18922 , \ILAB0102.net20974 , \ILAB0102.ILE0916.net2656 , 
    \ILAB0102.net18589 , \ILAB0102.net18184 , \ILAB0102.net25699 , \ILAB0102.net17636 , \ILAB0102.net17978 , \ILAB0102.net17977 , \ILAB0102.net17618 , \ILAB0102.net25223 , \ILAB0102.net17617 , \ILAB0102.ILE0809.net2656 , 
    \ILAB0102.net20588 , \ILAB0102.net17687 , \ILAB0102.net26349 , \ILAB0102.ILE1503.net0541 , \ILAB0102.ILE0405.net2656 , \ILAB0102.net17957 , \ILAB0102.net23109 , \ILAB0102.net23107 , \ILAB0102.net17799 , \ILAB0102.ILE1005.net2656 , 
    \net17226<1> , \net10348<0> , \net10387<1> , \ILAB0102.ILE1416.net01339 , \net10387<6> , \ILAB0102.net19372 , \net18532<1> , \ILAB0102.net17912 , \ILAB0102.net18814 , \ILAB0102.ILE1416.net2656 , 
    \ILAB0102.net24799 , \ILAB0102.net25224 , \ILAB0102.net22639 , \ILAB0102.net18002 , \ILAB0102.net18004 , \ILAB0102.ILE0808.net2656 , \ILAB0102.net25717 , \ILAB0102.net19552 , \ILAB0102.net18157 , \ILAB0102.net19507 , 
    \ILAB0102.net18067 , \ILAB0102.net25042 , \ILAB0102.ILE0406.net2656 , \net18572<1> , \ILAB0102.net18182 , \ILAB0102.ILE1506.net2656 , \ILAB0102.net22549 , \ILAB0102.net19102 , \ILAB0102.net25519 , \ILAB0102.ILE0513.net2656 , 
    \net10337<4> , \ILAB0102.net20407 , \ILAB0102.net19373 , \ILAB0102.net19417 , \ILAB0102.net18383 , \ILAB0102.ILE0409.net2656 , \ILAB0102.net22684 , \ILAB0102.net23602 , \ILAB0102.ILE0811.net2656 , \ILAB0102.net24637 , 
    \ILAB0102.net25942 , \ILAB0102.net24638 , \ILAB0102.net18517 , \ILAB0102.net18519 , \ILAB0102.ILE0908.net2656 , \ILAB0102.ILE0606.net2656 , \ILAB0102.net24660 , \ILAB0102.ILE0806.net2656 , \ILAB0102.net21784 , \ILAB0102.net21694 , 
    \ILAB0102.net21379 , \ILAB0102.net21692 , \ILAB0102.net18679 , \ILAB0102.net18949 , \ILAB0102.net18654 , \ILAB0102.ILE0812.net2656 , \ILAB0102.net21152 , \ILAB0102.ILE1306.net2656 , \ILAB0102.net26257 , \ILAB0102.ILE0506.net2656 , 
    \ILAB0102.net22028 , \ILAB0102.net19642 , \ILAB0102.ILE1516.net2656 , \net10356<0> , \net10419<0> , \net10419<5> , \ILAB0102.net19687 , \ILAB0102.ILE0616.net2656 , \ILAB0102.net23494 , \ILAB0102.ILE0814.net01345 , 
    \ILAB0102.ILE0814.net2656 , \ILAB0102.net23692 , \ILAB0102.net25312 , \ILAB0102.net21244 , \ILAB0102.net21690 , \ILAB0102.net19939 , \ILAB0102.net23872 , \ILAB0102.net19868 , \ILAB0102.net19867 , \ILAB0102.net19013 , 
    \ILAB0102.net19084 , \ILAB0102.ILE0412.net2656 , \ILAB0102.net19462 , \ILAB0102.net19463 , \ILAB0102.ILE0509.net2656 , \ILAB0102.net25494 , \ILAB0102.net23269 , \ILAB0102.ILE0914.net2656 , \ILAB0102.net21262 , \ILAB0102.net22144 , 
    \ILAB0102.net19804 , \ILAB0102.ILE0414.net2656 , \net10355<0> , \ILAB0102.net22406 , \ILAB0102.ILE0716.net01339 , \net10415<0> , \ILAB0102.net22388 , \net10415<6> , \ILAB0102.ILE0716.net2656 , \ILAB0102.ILE0613.net0562 , 
    \ILAB0102.ILE0613.net0558 , \ILAB0102.net19329 , \ILAB0102.ILE0613.net2656 , \net10337<3> , \net18548<1> , \ILAB0102.net19399 , \ILAB0102.net19622 , \ILAB0102.ILE0408.net2656 , \ILAB0102.net21062 , \ILAB0102.net19620 , 
    \ILAB0102.ILE0508.net2656 , \ILAB0102.net25764 , \ILAB0102.net21128 , \ILAB0102.net25627 , \net18564<1> , \ILAB0102.ILE1408.net2656 , \ILAB0102.ILE1508.net2656 , \ILAB0102.ILE0608.net2656 , \ILAB0102.net24116 , \ILAB0102.net19935 , 
    \ILAB0102.ILE0612.net2656 , \ILAB0102.ILE0514.net2656 , \ILAB0102.net19847 , \ILAB0102.ILE1414.net2656 , \ILAB0102.net21514 , \ILAB0102.net23874 , \ILAB0102.net21467 , \ILAB0102.ILE0411.net2656 , \ILAB0102.net24142 , \ILAB0102.net21488 , 
    \ILAB0102.net19913 , \ILAB0102.ILE0712.net2656 , \ILAB0102.net19976 , \ILAB0102.net21559 , \ILAB0102.net19959 , \ILAB0102.ILE0713.net2656 , \ILAB0102.net20831 , \ILAB0102.net20812 , \net17182<6> , \ILAB0102.ILE1403.net2656 , 
    \net18544<6> , \net17218<6> , \Fast_out_28<5> , \ILAB0102.ILE0503.net2656 , \net17222<3> , \net10430<6> , \ILAB0102.ILE0403.net2656 , \ILAB0102.ILE0204.net2656 , \ILAB0102.net20291 , \ILAB0102.net26168 , 
    \net17202<3> , \ILAB0102.ILE0903.net2656 , \ILAB0102.net26124 , \ILAB0102.ILE0803.net0558 , \ILAB0102.net20678 , \ILAB0102.ILE0803.net2656 , \ILAB0102.ILE0511.net2656 , \net18552<1> , \ILAB0102.net20434 , \ILAB0102.ILE1301.net01342 , 
    \ILAB0102.net20929 , \ILAB0102.net20704 , \net17214<5> , \ILAB0102.ILE0601.net01339 , \ILAB0102.net20612 , \ILAB0102.ILE0601.net2656 , \ILAB0102.ILE0601.net0541 , \ILAB0102.ILE0501.net01339 , \ILAB0102.net20634 , \ILAB0102.ILE0501.net2656 , 
    \net17206<5> , \ILAB0102.ILE0801.net01339 , \net17206<1> , \ILAB0102.ILE0801.net2656 , \ILAB0102.ILE0801.net0541 , \ILAB0102.ILE0401.net01339 , \ILAB0102.net20724 , \ILAB0102.ILE0401.net2656 , \ILAB0102.ILE1401.net01339 , \ILAB0102.ILE1501.net01339 , 
    \net17178<0> , \net17148<1> , \net17202<4> , \net17202<0> , \ILAB0102.ILE0901.net2656 , \net10391<1> , \net10391<0> , \net10391<5> , \ILAB0102.net23243 , \net10391<4> , 
    \ILAB0102.ILE1316.net2656 , \ILAB0102.net22207 , \ILAB0102.ILE0708.net2656 , \ILAB0102.net21352 , \ILAB0102.net21107 , \ILAB0102.net21109 , \ILAB0102.net25061 , \ILAB0102.net25628 , \ILAB0102.ILE1406.net2656 , \net10395<1> , 
    \ILAB0102.net24414 , \ILAB0102.ILE1216.net01339 , \ILAB0102.net21197 , \ILAB0102.ILE1216.net2656 , \ILAB0102.ILE1216.net0541 , \ILAB0102.ILE1312.net2656 , \ILAB0102.net21377 , \ILAB0102.ILE1212.net2656 , \ILAB0102.net21416 , \ILAB0102.net22657 , 
    \ILAB0102.net21667 , \ILAB0102.net24862 , \ILAB0102.ILE0611.net2656 , \ILAB0102.ILE0611.net0541 , \ILAB0102.ILE0711.net0562 , \ILAB0102.ILE0711.net2656 , \ILAB0102.net23017 , \net10399<0> , \net10403<1> , \ILAB0102.net24459 , 
    \net10403<2> , \net10403<3> , \ILAB0102.ILE1016.net2656 , \ILAB0102.ILE1608.net0562 , \ILAB0102.net22659 , \ILAB0102.net24863 , \ILAB0102.ILE1012.net2656 , \ILAB0102.net24504 , \net10399<3> , \net10399<5> , 
    \ILAB0102.ILE1116.net2656 , \ELLR15_28<3> , \ILAB0102.net22297 , \ILAB0102.ILE0216.net2656 , \ILAB0102.net24529 , \ILAB0102.net24484 , \ILAB0102.net22097 , \ILAB0102.net24482 , \ILAB0102.net22099 , \ILAB0102.net22189 , 
    \ILAB0102.ILE0815.net2656 , \ILAB0102.ILE0614.net2656 , \ILAB0102.net24527 , \ILAB0102.ILE0915.net2656 , \ILAB0102.net25537 , \ILAB0102.net23287 , \ILAB0102.net23989 , \ILAB0102.ILE0714.net2656 , \ILAB0102.ILE0714.net0541 , \ILAB0102.net24212 , 
    \ILAB0102.ILE0515.net2656 , \ILAB0102.ILE0515.net0541 , \net10431<1> , \net10431<3> , \ILAB0102.ILE0316.net01339 , \net10431<0> , \ILAB0102.ILE0316.net2656 , \ILAB0102.ILE0813.net2656 , \ILAB0102.ILE1011.net2656 , \net18536<0> , 
    \ILAB0102.ILE1415.net2656 , \ILAB0102.net25159 , \ILAB0102.ILE1104.net2656 , \ILAB0102.net23175 , \ILAB0102.ILE0213.net2656 , \ILAB0102.net23132 , \ILAB0102.ILE1004.net2656 , \ILAB0102.net23377 , \ILAB0102.net26100 , \ILAB0102.ILE0313.net2656 , 
    \ILAB0102.ILE0305.net2656 , \ILAB0102.net25898 , \ILAB0102.net23379 , \ILAB0102.ILE0311.net2656 , \ILAB0102.ILE1014.net2656 , \ILAB0102.ILE1014.net0541 , \ILAB0102.net24889 , \ILAB0102.net24754 , \ILAB0102.ILE0810.net2656 , \ILAB0102.ILE0810.net0541 , 
    \ILAB0102.net25314 , \ILAB0102.net24885 , \ILAB0102.ILE0910.net2656 , \ILAB0102.net26754 , \ILAB0102.ILE0203.net2656 , \ILAB0102.net24169 , \ILAB0102.net24124 , \ILAB0102.net23895 , \ILAB0102.ILE0410.net2656 , \ILAB0102.ILE0510.net0562 , 
    \ILAB0102.ILE0510.net0558 , \ILAB0102.ILE0510.net2656 , \ILAB0102.ILE0615.net2656 , \ILAB0102.net24079 , \ILAB0102.net24165 , \ILAB0102.ILE0610.net2656 , \ILAB0102.ILE0710.net2656 , \ILAB0102.ILE0715.net2656 , \ILAB0102.ILE0715.net0541 , \ILAB0102.ILE1315.net2656 , 
    \ILAB0102.ILE1215.net2656 , \ILAB0102.ILE1015.net2656 , \ILAB0102.ILE1115.net01345 , \ILAB0102.ILE1115.net2656 , \ELLR14_28<3> , \ILAB0102.ILE0215.net2656 , \ILAB0102.net25404 , \ILAB0102.ILE0906.net2656 , \ILAB0102.net24752 , \ILAB0102.ILE1210.net2656 , 
    \ILAB0102.ILE0315.net2656 , \ILAB0102.net24975 , \ILAB0102.ILE1010.net2656 , \ILAB0102.ILE0312.net2656 , \ILAB0102.ILE1110.net2656 , \ILAB0102.ILE0504.net2656 , \ILAB0102.net25629 , \ILAB0102.ILE1405.net2656 , \ILAB0102.ILE0904.net0541 , \ILAB0102.ILE1304.net2656 , 
    \ILAB0102.net25832 , \ILAB0102.ILE0807.net2656 , \ELLR9_28<5> , \ILAB0102.ILE0909.net2656 , \ILAB0102.ILE1604.net0558 , \ILAB0102.ILE1604.net0541 , \ILAB0102.ILE0905.net2656 , \ILAB0102.ILE0913.net2656 , \ILAB0102.ILE0804.net01345 , \ILAB0102.ILE0804.net2656 , 
    \ILAB0102.ILE1404.net2656 , \ILAB0102.ILE1507.net2656 , \ILAB0102.ILE1407.net2656 , \ILAB0102.net25830 , \ILAB0102.ILE1007.net2656 , \ILAB0102.ILE0310.net2656 , \ILAB0102.ILE0907.net2656 , \ILAB0102.ILE0604.net0562 , \ILAB0102.ILE0604.net2656 , \ILAB0102.ILE0413.net2656 , 
    \ILAB0102.net26689 , \ILAB0102.net26192 , \ILAB0102.net26599 , \ILAB0102.net26149 , \ILAB0102.ILE0802.net2656 , \ILAB0102.net26554 , \ILAB0102.ILE0902.net2656 , \ILAB0102.ILE0402.net2656 , \ILAB0102.ILE0502.net2656 , \net18588<0> , 
    \ILAB0102.net26509 , \net18588<1> , \ILAB0102.net26329 , \ILAB0102.ILE1402.net2656 , \ILAB0102.ILE1402.net0541 , \net18588<3> , \ILAB0102.ILE1502.net2656 , \ILAB0102.ILE0602.net2656 , \ILAB0102.ILE1602.net01339 , \net18588<6> , 
    \net18588<5> , \ILAB0102.ILE1602.net2656 , \ILAB0102.net26552 , \ILAB0102.ILE1302.net2656 , \ILAB0102.ILE1102.net2656 , \ILAB0102.ILE1102.net0541 , \ILAB0102.ILE0202.net2656 , \net16523<0> , \net16523<1> , \net16539<1> , 
    \net16578<1> , \ILAB0302.I5605.net21 , \ILAB0302.Clk_int<0> , \ILAB0302.net027160 , \ILAB0302.I5366.net70 , \net16372<0> , \ILAB0302.I5366.net0119 , \net16372<1> , \ILAB0302.I5366.net0110 , \ILAB0302.net15299<2> , 
    \ILAB0302.Clk_LAB<1> , \net16386<0> , \net16387<0> , \ILAB0302.net38580 , \ILAB0302.net20569 , \net11344<0> , \net11344<3> , \net11344<1> , \net11344<6> , \ILAB0302.ILE1601.net2656 , 
    \ILAB0302.ILE1501.net01339 , \ILAB0302.ILE1501.net2656 , \ILAB0302.ILE1501.net0541 , \ILAB0302.net26599 , \ILAB0302.net26149 , \net11189<6> , \ILAB0302.net26509 , \net11340<3> , \net11340<6> , \ILAB0402.I5366.net70 , 
    \ILAB0402.I5366.net0110 , \ILAB0402.net15299<2> , \ILAB0402.Clk_LAB<1> , \net16245<0> , \net16244<0> , \ILAB0402.net16736 , \ILAB0402.net37806 , \net16304<3> , \ILAB0402.net20587 , \net16328<1> , 
    \ILAB0402.net16719 , \ILAB0402.ILE0101.net2656 , \ILAB0402.net16961 , \net16324<4> , \net16324<5> , \net16324<1> , \ILAB0402.net16944 , \ILAB0402.ILE0201.net2656 , \net16308<3> , \net16248<1> , 
    \net16320<3> , \ILAB0402.ILE0301.net01339 , \net16320<2> , \ILAB0402.ILE0301.net2656 , \ILAB0402.net20651 , \net16312<3> , \net16244<1> , \ILAB0402.net20929 , \net16304<5> , \net16304<0> , 
    \ILAB0402.ILE0701.net0541 , \net16235<1> , \net16308<2> , \net16308<0> , \ILAB0402.net20612 , \ILAB0402.ILE0601.net0541 , \net16312<5> , \net16312<1> , \net16312<0> , \ILAB0402.ILE0501.net2656 , 
    \net16243<1> , \ILAB0402.ILE0401.net0562 , \ILAB0402.ILE0401.net0558 , \ILAB0402.ILE0401.net01342 , \ILAB0402.ILE0401.net2656 , \ILAB0402.net26419 , \net11247<1> , \ILAB0402.ILE0502.net0562 , \ILAB0402.ILE0502.net2656 , \ILAB0402.ILE0502.net0541 , 
    \ILAB0402.ILE0102.net01339 , \ILAB0402.net26775 , \ILAB0402.ILE0102.net2656 , \ILAB0402.ILE0102.net0541 , \ILAB0402.ILE0202.net2656 , \ILAB0402.ILE0202.net0541 , \ILAB0402.ILE0302.net2656 , \ILAB0103.I5605.net25 , \ILAB0103.Clk_int<1> , \ILAB0103.net027166 , 
    \ILAB0103.I5366.net66 , \ILAB0103.I5366.net0110 , \ILAB0103.net15299<2> , \ILAB0103.I5366.net0102 , \ILAB0103.net15299<0> , \ILAB0103.Clk_LAB<1> , \ILAB0103.Clk_LAB<3> , \ILAB0103.net15476 , \ILAB0103.net26501 , \ILAB0103.net20561 , 
    \ILAB0103.net38382 , \ILAB0103.net37923 , \ILAB0103.net37740 , \ILAB0103.net39618 , \ILAB0103.net22946 , \ILAB0103.net38496 , \ILAB0103.net22856 , \ILAB0103.net37425 , \ILAB0103.net39588 , \ILAB0103.net39060 , 
    \net18735<3> , \ILAB0103.net20884 , \ILAB0103.net15502 , \ILAB0103.net15504 , \ILAB0103.ILE1201.net2656 , \ILAB0103.net16114 , \ILAB0103.net25609 , \net11483<6> , \Fast_out_29<4> , \ILAB0103.ILE0404.net2656 , 
    \ILAB0103.net17734 , \ILAB0103.net26574 , \ILAB0103.net26573 , \ILAB0103.net15594 , \ILAB0103.ILE1203.net2656 , \ILAB0103.net20299 , \ILAB0103.net20497 , \ILAB0103.net26438 , \ILAB0103.net26437 , \ILAB0103.net16924 , 
    \ILAB0103.net15709 , \ILAB0103.net20344 , \ILAB0103.net15684 , \ILAB0103.ILE0703.net2656 , \ILAB0103.net17374 , \ILAB0103.net25989 , \ILAB0103.net15799 , \ILAB0103.net15844 , \ILAB0103.ILE0605.net2656 , \ILAB0103.ILE0705.net2656 , 
    \ILAB0103.net20452 , \ILAB0103.net23134 , \ILAB0103.net25114 , \ILAB0103.net25112 , \ILAB0103.ILE0704.net2656 , \net18731<1> , \ILAB0103.net16556 , \ILAB0103.ILE1001.net2656 , \ILAB0103.ILE1101.net01345 , \ILAB0103.net16583 , 
    \ILAB0103.ILE1101.net2656 , \net11495<6> , \Fast_out_29<7> , \ILAB0103.net24997 , \ILAB0103.net26664 , \ILAB0103.ILE1103.net2656 , \ILAB0103.ILE0201.net01339 , \ILAB0103.net20614 , \ILAB0103.net17865 , \ILAB0103.ILE0201.net2656 , 
    \ILAB0103.net25584 , \ILAB0103.ILE0805.net2656 , \ILAB0103.net26618 , \ILAB0103.net17394 , \ILAB0103.ILE1003.net2656 , \ILAB0103.net20606 , \ILAB0103.net20524 , \ILAB0103.ILE0301.net2656 , \ILAB0103.net26752 , \ILAB0103.net20632 , 
    \ILAB0103.net26259 , \ILAB0103.net26276 , \ILAB0103.net20633 , \ILAB0103.net20162 , \Fast_out_29<5> , \ILAB0103.ILE0503.net2656 , \ILAB0103.ILE0503.net0541 , \ILAB0103.net26214 , \net11487<6> , \ILAB0103.ILE0403.net2656 , 
    \ILAB0103.net26168 , \ILAB0103.net20274 , \ILAB0103.ILE0903.net2656 , \ILAB0103.net20678 , \ILAB0103.net20454 , \ILAB0103.ILE1301.net2656 , \ILAB0103.net20929 , \ILAB0103.ILE0701.net01345 , \ILAB0103.ILE0701.net01339 , \ILAB0103.net20522 , 
    \ILAB0103.ILE0701.net2656 , \ILAB0103.net20612 , \ILAB0103.ILE0601.net2656 , \ILAB0103.net20655 , \ILAB0103.ILE0501.net2656 , \ILAB0103.net20679 , \ILAB0103.ILE0801.net2656 , \ILAB0103.ILE0401.net01339 , \ILAB0103.ILE0401.net2656 , \ILAB0103.ILE0401.net0541 , 
    \ILAB0103.ILE0901.net2656 , \net11487<3> , \ILAB0103.net25654 , \ILAB0103.ILE1204.net2656 , \ILAB0103.net23132 , \ILAB0103.ILE1004.net2656 , \ILAB0103.ILE0303.net2656 , \ILAB0103.net24999 , \ILAB0103.ILE0504.net2656 , \ILAB0103.ILE0904.net2656 , 
    \ILAB0103.ILE0505.net2656 , \ILAB0103.ILE0804.net2656 , \ILAB0103.ILE0604.net2656 , \ILAB0103.net26644 , \ILAB0103.net26192 , \ILAB0103.net26149 , \ILAB0103.net26194 , \ILAB0103.ILE0802.net2656 , \ILAB0103.net26554 , \ILAB0103.ILE0902.net2656 , 
    \ILAB0103.net26464 , \ILAB0103.ILE0402.net0562 , \ILAB0103.ILE0402.net0558 , \ILAB0103.ILE0402.net2656 , \ILAB0103.ILE0502.net2656 , \ILAB0103.net26329 , \ILAB0103.ILE0602.net2656 , \ILAB0103.ILE0602.net0541 , \ILAB0103.ILE0702.net2656 , \ILAB0103.ILE1602.net0560 , 
    \ILAB0103.ILE1302.net2656 , \ILAB0103.ILE1202.net2656 , \ILAB0103.ILE1002.net0541 , \ILAB0103.ILE1102.net2656 , \ILAB0103.ILE0302.net2656 , \Fast_in_32<7> , \ILAB0401.I5605.net25 , \ILAB0401.Clk_int<1> , \ILAB0401.I5605.net29 , \ILAB0401.Clk_int<3> , 
    \ILAB0401.I5605.net33 , \ILAB0401.Clk_int<2> , \ILAB0401.net027166 , \ILAB0401.net27188 , \ILAB0401.net015238 , \ILAB0401.I5366.net64 , \ILAB0401.I5366.net0114 , \ILAB0401.net15299<3> , \ILAB0401.I5366.net0110 , \ILAB0401.net15299<2> , 
    \ILAB0401.I5366.net0106 , \ILAB0401.net15299<1> , \ILAB0401.I5366.net0102 , \ILAB0401.net15299<0> , \ILAB0401.Clk_LAB<0> , \ILAB0401.Clk_LAB<1> , \ILAB0401.Clk_LAB<2> , \ILAB0401.Clk_LAB<3> , \ILAB0401.net27305 , \ILAB0401.net27353 , 
    \ILAB0401.net21911 , \ILAB0401.net15656 , \ILAB0401.net17212 , \ILAB0401.net21037 , \ILAB0401.net15637 , \ILAB0401.net24322 , \ILAB0401.net16312 , \ILAB0401.net17464 , \ILAB0401.net19309 , \ILAB0401.net19057 , 
    \ILAB0401.net17014 , \ILAB0401.ILE0516.net2656 , \ILAB0401.ILE0416.net01342 , \ILAB0401.net19238 , \ILAB0401.ILE0416.net2656 , \ILAB0401.net21604 , \ILAB0401.ILE0816.net01339 , \ILAB0401.ILE0816.net01342 , \ILAB0401.ILE0916.net01345 , \ILAB0401.ILE0916.net01339 , 
    \ILAB0401.net18922 , \ILAB0401.net17636 , \ILAB0401.net17977 , \ILAB0401.net18311 , \ILAB0401.net18315 , \ILAB0401.net19076 , \ILAB0401.net23917 , \ILAB0401.net18293 , \ILAB0401.net20363 , \ILAB0401.net19102 , 
    \ILAB0401.net25519 , \ILAB0401.net18319 , \ILAB0401.net19354 , \ILAB0401.net19350 , \ILAB0401.ILE0513.net2656 , \ILAB0401.ILE0513.net0541 , \ILAB0401.net23044 , \ILAB0401.net22684 , \ILAB0401.net18992 , \ILAB0401.ILE0811.net01345 , 
    \ILAB0401.net18472 , \ILAB0401.net18499 , \ILAB0401.ILE0811.net2656 , \ILAB0401.net21694 , \ILAB0401.net18653 , \ILAB0401.net18677 , \ILAB0401.net18679 , \ILAB0401.net18949 , \ILAB0401.ILE0812.net2656 , \ILAB0401.net23964 , 
    \ILAB0401.ILE0616.net0558 , \ILAB0401.ILE0616.net2656 , \ILAB0401.net23494 , \ILAB0401.net22524 , \ILAB0401.net22541 , \ILAB0401.net18904 , \ILAB0401.net19174 , \ILAB0401.ILE0814.net2656 , \ILAB0401.ILE0814.net0541 , \ILAB0401.net23711 , 
    \ILAB0401.net18968 , \ILAB0401.net25312 , \ILAB0401.net18924 , \ILAB0401.ILE0912.net2656 , \ILAB0401.net25313 , \ILAB0401.net23042 , \ILAB0401.net22680 , \ILAB0401.ILE0911.net2656 , \ILAB0401.ILE0911.net0541 , \ILAB0401.net19939 , 
    \ILAB0401.net19714 , \ILAB0401.net19867 , \ILAB0401.net19084 , \ILAB0401.ILE0412.net2656 , \ILAB0401.ILE0512.net2656 , \ILAB0401.net25494 , \ILAB0401.net23269 , \ILAB0401.ILE0914.net2656 , \ILAB0401.net22414 , \ILAB0401.net22144 , 
    \ILAB0401.net19802 , \ILAB0401.net26078 , \net16275<6> , \ILAB0401.net19804 , \ILAB0401.ILE0414.net2656 , \ILAB0401.ILE0716.net01339 , \ILAB0401.net22388 , \ILAB0401.ILE0716.net2656 , \ILAB0401.net19346 , \ILAB0401.net19706 , 
    \ILAB0401.net19328 , \ILAB0401.net21424 , \ILAB0401.ILE0613.net2656 , \ILAB0401.ILE0613.net0541 , \ILAB0401.ILE0612.net01342 , \ILAB0401.ILE0612.net2656 , \ILAB0401.net22412 , \ILAB0401.ILE0514.net2656 , \ILAB0401.net21514 , \ILAB0401.net21487 , 
    \ILAB0401.net19913 , \ILAB0401.net24143 , \ILAB0401.net19914 , \ILAB0401.ILE0712.net2656 , \ILAB0401.net19976 , \ILAB0401.ILE0713.net0560 , \ILAB0401.net21559 , \ILAB0401.ILE0713.net2656 , \ILAB0401.ILE1601.net01345 , \ILAB0401.ILE1616.net01345 , 
    \ILAB0401.net22657 , \ILAB0401.net21669 , \ILAB0401.ILE1013.net2656 , \ILAB0401.ILE0611.net2656 , \ILAB0401.ILE0711.net0558 , \ILAB0401.ILE0711.net2656 , \ILAB0401.ILE1016.net01345 , \ILAB0401.ILE1016.net01342 , \ILAB0401.ILE1012.net2656 , \net16267<3> , 
    \ILAB0401.net24549 , \ILAB0401.ILE0116.net01339 , \ILAB0401.net23648 , \ILAB0401.net21892 , \ILAB0401.ILE0116.net2656 , \net16283<3> , \ILAB0401.net25267 , \ILAB0401.net23197 , \ILAB0401.ILE0216.net2656 , \ILAB0401.net22189 , 
    \ILAB0401.net22119 , \ILAB0401.ILE0614.net2656 , \ILAB0401.ILE0614.net0541 , \net16279<6> , \net16279<3> , \ILAB0401.ILE0113.net01339 , \ILAB0401.net22253 , \ILAB0401.net23177 , \net16279<1> , \ILAB0401.net22254 , 
    \ILAB0401.ILE0113.net2656 , \ILAB0401.ILE0113.net0541 , \ILAB0401.net25537 , \ILAB0401.net24930 , \ILAB0401.ILE0212.net2656 , \ILAB0401.net22365 , \net16271<6> , \ILAB0401.ILE0415.net2656 , \ILAB0401.ILE0714.net01339 , \ILAB0401.ILE0714.net0541 , 
    \ILAB0401.ILE0515.net2656 , \ILAB0401.net23801 , \ILAB0401.ILE0316.net01342 , \ILAB0401.net24907 , \ILAB0401.ILE0316.net2656 , \ILAB0401.ILE0316.net0541 , \ILAB0401.ILE0813.net01339 , \ILAB0401.ILE0813.net2656 , \ILAB0401.ILE1011.net2656 , \ILAB0401.net26102 , 
    \ILAB0401.net23175 , \ILAB0401.ILE0213.net2656 , \ILAB0401.net23396 , \ILAB0401.net23377 , \ILAB0401.net24908 , \ILAB0401.net23153 , \ILAB0401.net23154 , \ILAB0401.ILE0313.net2656 , \ILAB0401.ILE1014.net2656 , \ILAB0401.net24979 , 
    \ILAB0401.net24889 , \ILAB0401.net23717 , \ILAB0401.net23719 , \ILAB0401.ILE0810.net0541 , \ILAB0401.ILE0114.net2656 , \ILAB0401.net24977 , \ILAB0401.net24885 , \ILAB0401.ILE0910.net2656 , \ILAB0401.ILE0214.net01339 , \ILAB0401.ILE0214.net2656 , 
    \ILAB0401.net23784 , \ILAB0401.ILE0314.net2656 , \ILAB0401.ILE0615.net2656 , \ILAB0401.ILE0710.net2656 , \ILAB0401.ILE0710.net0541 , \ILAB0401.ILE0715.net01339 , \ILAB0401.ILE0715.net2656 , \net16271<1> , \ILAB0401.ILE0115.net2656 , \ILAB0401.ILE0215.net2656 , 
    \ILAB0401.net24752 , \ILAB0401.ILE0315.net2656 , \ILAB0401.ILE0315.net0541 , \ILAB0401.ILE1010.net01342 , \ILAB0401.ILE1010.net2656 , \ILAB0401.ILE0312.net2656 , \ILAB0401.ILE0312.net0541 , \ILAB0401.ILE0913.net2656 , \ILAB0401.ILE0413.net01345 , \ILAB0401.ILE0413.net2656 , 
    \ILAB0301.I5605.net29 , \ILAB0301.Clk_int<3> , \ILAB0301.net015234 , \ILAB0301.I5366.net0122 , \ILAB0301.net22766 , \ILAB0301.net19354 , \net16377<4> , \ILAB0301.net18364 , \ILAB0301.net21424 , \net16430<1> , 
    \ILAB1001.I5605.net21 , \ILAB1001.Clk_int<0> , \ILAB1001.I5605.net25 , \ILAB1001.Clk_int<1> , \ILAB1001.net027160 , \ILAB1001.net027166 , \ILAB1001.I5366.net68 , \ILAB1001.I5366.net0122 , \ILAB1001.I5366.net0119 , \ILAB1001.I5366.net0106 , 
    \ILAB1001.net15299<1> , \ILAB1001.Clk_LAB<2> , \ILAB1001.net20561 , \ILAB1001.net27361 , \ILAB1001.net25762 , \ILAB1001.net21127 , \ILAB1001.net24007 , \ILAB1001.net26302 , \ILAB1001.net20002 , \ILAB1001.ILE1403.net2656 , 
    \ILAB1001.ILE1410.net2656 , \ILAB1001.ILE1610.net0562 , \ILAB0101.I5366.net64 , \ILAB0101.I5366.net0114 , \ILAB0101.net15299<3> , \ILAB0101.Clk_LAB<0> , \ILAB0101.net27295 , \ILAB0101.net27297 , \ILAB0101.ILE0416.net01342 , \ILAB0101.ILE0916.net2656 , 
    \ILAB0101.ILE0916.net0541 , \net17132<4> , \ILAB0101.ILE1516.net01345 , \ILAB0101.ILE1516.net01342 , \ILAB0101.ILE1513.net2656 , \ILAB0101.ILE1613.net0562 , \ILAB0101.net23756 , \ILAB0101.ILE0216.net01339 , \net18389<6> , \ILAB0101.ILE0215.net0541 , 
    \ILAB0201.I5366.net64 , \ILAB0201.I5366.net0114 , \ILAB0201.net15299<3> , \ILAB0201.Clk_LAB<0> , \net18362<1> , \ILAB0201.net27303 , \ILAB0201.net19354 , \ILAB0201.net18364 , \ILAB0201.net21424 , \ILAB0201.ILE0316.net01345 , 
    \ILAB0201.ILE0316.net01339 , \ILAB0201.net25897 , \ILAB0201.net23154 , \ILAB0201.ILE0313.net2656 , \ILAB0201.net23807 , \ILAB0201.ILE0314.net2656 , \ILAB0202.I5366.net68 , \ILAB0202.I5366.net70 , \ILAB0202.I5366.net0110 , \ILAB0202.net15299<2> , 
    \ILAB0202.I5366.net0106 , \ILAB0202.net15299<1> , \ILAB0202.Clk_LAB<1> , \ILAB0202.Clk_LAB<2> , \ILAB0202.net23216 , \ILAB0202.net40041 , \ILAB0202.net21911 , \ILAB0202.net38625 , \ILAB0202.net19732 , \ILAB0202.net16718 , 
    \ILAB0202.net22837 , \ILAB0202.ILE0106.net01339 , \ILAB0202.ILE0105.net2656 , \ILAB0202.ILE0205.net2656 , \ILAB0202.ILE0103.net01345 , \ILAB0202.ILE0103.net01342 , \ILAB0202.ILE0103.net2656 , \ILAB0202.ILE0108.net01339 , \ILAB0202.net26599 , \ILAB0202.net26149 , 
    \ILAB0202.net26509 , \ILAB0202.net26822 , \ILAB0202.ILE0202.net2656 , \ILAB0202.ILE0302.net2656 , \IIO31.net728 , \IIO12.I7.net197 , \IIO12.I6.net197 , \IIO12.I5.net197 , \IIO12.I4.net197 , \IIO12.I3.net197 , 
    \IIO12.I2.net197 , \IIO12.I1.net197 , \IIO12.I0.net197 , \IIO33.I6.net0153 , \IIO33.I6.net209 , \IIO33.I5.net0151 , \IIO33.I5.net0153 , \IIO33.I5.net209 , \IIO33.I4.net0153 , \IIO33.I4.net209 , 
    \IIO33.I3.net0153 , \IIO33.I3.net209 , \IIO33.I2.net0151 , \IIO33.I2.net0153 , \IIO33.I2.net209 , \IIO33.I1.net0153 , \IIO33.I1.net209 , \IIO33.I0.net0151 , \IIO33.I0.net0153 , \IIO33.I0.net209 , 
    \IIO13.I5.net197 , \IIO13.I4.net197 , \IIO13.I3.net197 , \IIO13.I2.net197 , \IIO13.I1.net197 , \IIO13.I0.net197 , \IIO10.I7.net197 , \IIO10.I6.net197 , \IIO10.I5.net197 , \IIO10.I4.net197 , 
    \IIO10.I3.net197 , \IIO10.I2.net197 , \IIO10.I1.net197 , \IIO11.I7.net197 , \IIO11.I6.net197 , \IIO11.I5.net197 , \IIO11.I4.net197 , \IIO11.I3.net197 , \IIO11.I2.net197 , \IIO11.I1.net197 , 
    \IIO11.I0.net197 ,
    GND, VDD;
  assign GND = 1'b0;
  assign VDD = 1'b1;

  //initial $sdf_annotate("C:/Users/Admin-PC/Desktop/sny/adc1_plasvet/adc_045/adc045_wrap.STA.reports/adc045_wrap.routed.sdf");

  xci2_ib XC_BUF_cs ( .a(cs), .x(\IIO33.I0.net209 ));
  xci2_ib XC_BUF_dout ( .a(dout), .x(\IIO33.I1.net209 ));
  xci2_ib XC_BUF_drdy ( .a(drdy), .x(\IIO33.I2.net209 ));
  xci2_ib XC_BUF_hard_start ( .a(hard_start), .x(\IIO33.I3.net209 ));
  xci2_ib XC_BUF_hard_wreg ( .a(hard_wreg), .x(\IIO33.I4.net209 ));
  xci2_ib XC_BUF_rst_l ( .a(rst_l), .x(\IIO33.I5.net209 ));
  xci2_ib XC_BUF_rst_l_adc ( .a(rst_l_adc), .x(\IIO33.I6.net209 ));
  xci2_ob XC_BUF_din ( .a(\IIO10.I1.net197 ), .x(din));
  xci2_ob XC_BUF_nRST ( .a(\IIO10.I2.net197 ), .x(nRST));
  xci2_ob XC_BUF_ready_sample ( .a(\IIO10.I3.net197 ), .x(ready_sample));
  xci2_ob XC_BUF_sclk ( .a(\IIO10.I4.net197 ), .x(sclk));
  xci2_ob XC_BUF_start ( .a(\IIO10.I5.net197 ), .x(start));
  xci2_ob \XC_BUF_adc045_data[0]  ( .a(\IIO10.I6.net197 ), .x(adc045_data[0]));
  xci2_ob \XC_BUF_adc045_data[10]  ( .a(\IIO10.I7.net197 ), .x(adc045_data[10]));
  xci2_ob \XC_BUF_adc045_data[11]  ( .a(\IIO11.I0.net197 ), .x(adc045_data[11]));
  xci2_ob \XC_BUF_adc045_data[12]  ( .a(\IIO11.I1.net197 ), .x(adc045_data[12]));
  xci2_ob \XC_BUF_adc045_data[13]  ( .a(\IIO11.I2.net197 ), .x(adc045_data[13]));
  xci2_ob \XC_BUF_adc045_data[14]  ( .a(\IIO11.I3.net197 ), .x(adc045_data[14]));
  xci2_ob \XC_BUF_adc045_data[15]  ( .a(\IIO11.I4.net197 ), .x(adc045_data[15]));
  xci2_ob \XC_BUF_adc045_data[16]  ( .a(\IIO11.I5.net197 ), .x(adc045_data[16]));
  xci2_ob \XC_BUF_adc045_data[17]  ( .a(\IIO11.I6.net197 ), .x(adc045_data[17]));
  xci2_ob \XC_BUF_adc045_data[18]  ( .a(\IIO11.I7.net197 ), .x(adc045_data[18]));
  xci2_ob \XC_BUF_adc045_data[19]  ( .a(\IIO12.I0.net197 ), .x(adc045_data[19]));
  xci2_ob \XC_BUF_adc045_data[1]  ( .a(\IIO12.I1.net197 ), .x(adc045_data[1]));
  xci2_ob \XC_BUF_adc045_data[20]  ( .a(\IIO12.I2.net197 ), .x(adc045_data[20]));
  xci2_ob \XC_BUF_adc045_data[21]  ( .a(\IIO12.I3.net197 ), .x(adc045_data[21]));
  xci2_ob \XC_BUF_adc045_data[22]  ( .a(\IIO12.I4.net197 ), .x(adc045_data[22]));
  xci2_ob \XC_BUF_adc045_data[23]  ( .a(\IIO12.I5.net197 ), .x(adc045_data[23]));
  xci2_ob \XC_BUF_adc045_data[2]  ( .a(\IIO12.I6.net197 ), .x(adc045_data[2]));
  xci2_ob \XC_BUF_adc045_data[3]  ( .a(\IIO12.I7.net197 ), .x(adc045_data[3]));
  xci2_ob \XC_BUF_adc045_data[4]  ( .a(\IIO13.I0.net197 ), .x(adc045_data[4]));
  xci2_ob \XC_BUF_adc045_data[5]  ( .a(\IIO13.I1.net197 ), .x(adc045_data[5]));
  xci2_ob \XC_BUF_adc045_data[6]  ( .a(\IIO13.I2.net197 ), .x(adc045_data[6]));
  xci2_ob \XC_BUF_adc045_data[7]  ( .a(\IIO13.I3.net197 ), .x(adc045_data[7]));
  xci2_ob \XC_BUF_adc045_data[8]  ( .a(\IIO13.I4.net197 ), .x(adc045_data[8]));
  xci2_ob \XC_BUF_adc045_data[9]  ( .a(\IIO13.I5.net197 ), .x(adc045_data[9]));
  xci2_ib_gclk XC_BUF_clk ( .a(clk), .x(\Fast_in_32<7> ));
  xci2_inv _184_ ( .a(\ILAB1001.net26302 ), .y(\ILAB1001.ILE1403.net2656 ));
  xci2_and2ft _185_ ( .a(\ILAB0102.net15864 ), .b(\ILAB0102.net15863 ), .y(\ILAB0202.ILE0205.net2656 ));
  xci2_and3ftt _186_ ( .a(\ILAB0101.ILE1613.net0562 ), .b(\ILAB0101.ILE1516.net01345 ), .c(\net17132<4> ), .y(\ILAB0101.ILE1513.net2656 ));
  xci2_nor2 _187_ ( .a(\ILAB0401.net23154 ), .b(\net16324<1> ), .y(\ILAB0401.ILE0314.net2656 ));
  xci2_and2ft _188_ ( .a(\ILAB0401.ILE0413.net01345 ), .b(\ILAB0401.net18319 ), .y(\ILAB0401.ILE0413.net2656 ));
  xci2_and3fft _189_ ( .a(\ILAB0401.net24907 ), .b(\ILAB0401.net26102 ), .c(\ILAB0401.net24549 ), .y(\ILAB0401.ILE0215.net2656 ));
  xci2_or3 _190_ ( .a(\ILAB0401.net19309 ), .b(\net11247<1> ), .c(\ILAB0402.net26419 ), .y(\ILAB0402.ILE0302.net2656 ));
  xci2_nor2ft _191_ ( .a(\ILAB0202.Clk_LAB<1> ), .b(\net18588<6> ), .y(\ILAB0202.ILE0202.net2656 ));
  xci2_or3fft _192_ ( .a(\ILAB0202.Clk_LAB<2> ), .b(\ILAB0202.Clk_LAB<1> ), .c(\net18588<6> ), .y(\ILAB0202.ILE0302.net2656 ));
  xci2_or2 _193_ ( .a(\ILAB0102.ILE1401.net01339 ), .b(\ILAB0102.Clk_LAB<2> ), .y(\ILAB0102.ILE1402.net2656 ));
  xci2_or2 _193__1 ( .a(\ILAB0102.ILE1401.net01339 ), .b(\ILAB0102.Clk_LAB<2> ), .y(\ILAB0102.ILE1402.net0541 ));
  xci2_nor3 _194_ ( .a(\ILAB0202.ILE0103.net01345 ), .b(\net18389<6> ), .c(\ILAB0102.Clk_LAB<2> ), .y(\ILAB0102.ILE1403.net2656 ));
  xci2_oa21ttf _195_ ( .a(\ILAB0202.ILE0103.net01345 ), .b(\ILAB0202.ILE0103.net01342 ), .c(\ILAB0202.net16718 ), .y(\ILAB0202.ILE0103.net2656 ));
  xci2_aoi21 _196_ ( .a(\ILAB0102.net26349 ), .b(\ILAB0102.net15482 ), .c(\ILAB0102.net20857 ), .y(\ILAB0102.ILE1503.net0541 ));
  xci2_oai21 _197_ ( .a(\net18389<6> ), .b(\net18588<3> ), .c(\ILAB0102.ILE1602.net01339 ), .y(\ILAB0102.ILE1602.net2656 ));
  xci2_ao21ftt _198_ ( .a(\net18588<0> ), .b(\ILAB0102.ILE1303.net0560 ), .c(\net18389<6> ), .y(\ILAB0102.ILE1303.net2656 ));
  xci2_nand2 _199_ ( .a(\ILAB0102.net15754 ), .b(\ILAB0101.ILE1516.net01342 ), .y(\ILAB0102.ILE1304.net2656 ));
  xci2_and3 _200_ ( .a(\ILAB0102.net26349 ), .b(\ILAB0102.net16654 ), .c(\ILAB0102.net25159 ), .y(\ILAB0102.ILE0905.net2656 ));
  xci2_ao21 _201_ ( .a(\ILAB0102.net24660 ), .b(\ILAB0102.net17799 ), .c(\ILAB0102.net25404 ), .y(\ILAB0102.ILE0906.net2656 ));
  xci2_and3 _202_ ( .a(\ILAB0102.net23692 ), .b(\ILAB0102.net25312 ), .c(\ILAB0102.net18922 ), .y(\ILAB0102.ILE0913.net2656 ));
  xci2_ao21 _203_ ( .a(\ILAB0102.net23494 ), .b(\ILAB0102.net22657 ), .c(\ILAB0102.net25494 ), .y(\ILAB0102.ILE0914.net2656 ));
  xci2_and3 _204_ ( .a(\ILAB0102.ILE1115.net01345 ), .b(\ILAB0102.net23017 ), .c(\net10391<0> ), .y(\ILAB0102.ILE1115.net2656 ));
  xci2_ao21 _205_ ( .a(\ILAB0103.ILE1101.net01345 ), .b(\ILAB0102.net19372 ), .c(\ILAB0102.net24504 ), .y(\ILAB0102.ILE1116.net2656 ));
  xci2_and3 _206_ ( .a(\ILAB0103.ILE1101.net01345 ), .b(\net10399<3> ), .c(\net10399<0> ), .y(\ILAB0103.ILE1101.net2656 ));
  xci2_ao21 _207_ ( .a(\net10395<1> ), .b(\net10387<6> ), .c(\ILAB0103.net20884 ), .y(\ILAB0103.ILE1201.net2656 ));
  xci2_and3 _208_ ( .a(\net10395<1> ), .b(\net10407<0> ), .c(\net10407<2> ), .y(\ILAB0103.ILE0901.net2656 ));
  xci2_ao21 _209_ ( .a(\net10411<1> ), .b(\net10403<3> ), .c(\ILAB0103.net20929 ), .y(\ILAB0103.ILE0801.net2656 ));
  xci2_and3 _210_ ( .a(\ILAB0103.net20678 ), .b(\net10403<1> ), .c(\net10407<2> ), .y(\ILAB0103.ILE1001.net2656 ));
  xci2_ao21 _211_ ( .a(\ILAB0102.net24459 ), .b(\net10403<3> ), .c(\net10403<2> ), .y(\ILAB0102.ILE1016.net2656 ));
  xci2_and3 _212_ ( .a(\ILAB0102.net24482 ), .b(\net10407<0> ), .c(\ILAB0102.net18922 ), .y(\ILAB0102.ILE0915.net2656 ));
  xci2_ao21 _213_ ( .a(\net10407<1> ), .b(\net10403<3> ), .c(\ILAB0102.net22164 ), .y(\ILAB0102.ILE0916.net2656 ));
  xci2_and3 _214_ ( .a(\net10407<1> ), .b(\ILAB0102.net23017 ), .c(\ILAB0102.net18878 ), .y(\ILAB0102.ILE0816.net2656 ));
  xci2_ao21 _215_ ( .a(\ILAB0102.net24529 ), .b(\ILAB0102.Clk_LAB<1> ), .c(\ILAB0102.net18652 ), .y(\ILAB0102.ILE0815.net2656 ));
  xci2_and3 _216_ ( .a(\ILAB0102.ILE0814.net01345 ), .b(\ILAB0102.net23017 ), .c(\ILAB0102.net21379 ), .y(\ILAB0102.ILE0814.net2656 ));
  xci2_ao21 _217_ ( .a(\ILAB0102.net17636 ), .b(\ILAB0102.Clk_LAB<1> ), .c(\ILAB0102.net23602 ), .y(\ILAB0102.ILE0811.net2656 ));
  xci2_and3 _218_ ( .a(\ILAB0102.net17978 ), .b(\ILAB0102.net17167 ), .c(\ILAB0102.net17347 ), .y(\ILAB0102.ILE0809.net2656 ));
  xci2_ao21 _219_ ( .a(\ILAB0102.net25832 ), .b(\ILAB0102.net17957 ), .c(\ILAB0102.net25223 ), .y(\ILAB0102.ILE0907.net2656 ));
  xci2_and3 _220_ ( .a(\ILAB0102.net23107 ), .b(\ILAB0102.net16652 ), .c(\ILAB0102.net25159 ), .y(\ILAB0102.ILE1104.net2656 ));
  xci2_ao21 _221_ ( .a(\ILAB0102.net26662 ), .b(\ILAB0102.net20029 ), .c(\net17194<6> ), .y(\ILAB0102.ILE1103.net2656 ));
  xci2_and3 _222_ ( .a(\ILAB0102.ILE1003.net0562 ), .b(\ILAB0102.net16654 ), .c(\ILAB0102.net25159 ), .y(\ILAB0102.ILE1003.net2656 ));
  xci2_ao21 _223_ ( .a(\ILAB0102.net26168 ), .b(\ILAB0102.net20029 ), .c(\ILAB0102.net17419 ), .y(\ILAB0102.ILE0903.net2656 ));
  xci2_and3 _224_ ( .a(\ILAB0102.net26168 ), .b(\ILAB0102.net16654 ), .c(\ILAB0102.net25114 ), .y(\ILAB0102.ILE0904.net0541 ));
  xci2_ao21 _225_ ( .a(\ILAB0102.net20340 ), .b(\ILAB0102.net20029 ), .c(\ILAB0102.ILE0803.net0558 ), .y(\ILAB0102.ILE0803.net2656 ));
  xci2_and3 _226_ ( .a(\ILAB0102.ILE0804.net01345 ), .b(\ILAB0102.net16654 ), .c(\ILAB0102.net25114 ), .y(\ILAB0102.ILE0804.net2656 ));
  xci2_ao21 _227_ ( .a(\ILAB0102.net17959 ), .b(\ILAB0102.net20029 ), .c(\ILAB0102.net25584 ), .y(\ILAB0102.ILE0805.net2656 ));
  xci2_and3 _228_ ( .a(\ILAB0102.net17214 ), .b(\ILAB0102.net16654 ), .c(\ILAB0102.net17347 ), .y(\ILAB0102.ILE0807.net2656 ));
  xci2_ao21 _229_ ( .a(\ILAB0102.net24799 ), .b(\ILAB0102.net17799 ), .c(\ILAB0102.net25224 ), .y(\ILAB0102.ILE0808.net2656 ));
  xci2_and3 _230_ ( .a(\ILAB0102.net24799 ), .b(\ILAB0102.net24638 ), .c(\ILAB0102.net25159 ), .y(\ILAB0102.ILE0908.net2656 ));
  xci2_ao21 _231_ ( .a(\ILAB0102.net25942 ), .b(\ILAB0102.net25807 ), .c(\ILAB0102.net18519 ), .y(\ILAB0102.ILE0909.net2656 ));
  xci2_and3 _232_ ( .a(\ILAB0102.net24885 ), .b(\ILAB0102.net18202 ), .c(\ILAB0102.net16222 ), .y(\ILAB0102.ILE1010.net2656 ));
  xci2_ao21 _233_ ( .a(\ILAB0102.net24754 ), .b(\ILAB0102.net19507 ), .c(\ILAB0102.net24975 ), .y(\ILAB0102.ILE1110.net2656 ));
  xci2_ao21 _234_ ( .a(\ILAB0202.net26822 ), .b(\ILAB0202.net22837 ), .c(\net18576<3> ), .y(\ILAB0202.ILE0105.net2656 ));
  xci2_nand3ftt _235_ ( .a(\ILAB0102.ILE1604.net0558 ), .b(\net18588<1> ), .c(\net18584<2> ), .y(\ILAB0102.ILE1504.net2656 ));
  xci2_ao21ttf _236_ ( .a(\ILAB0102.net17032 ), .b(\ILAB0202.net19732 ), .c(\ILAB0102.net16177 ), .y(\ILAB0102.ILE1507.net2656 ));
  xci2_ao21 _237_ ( .a(\net18572<1> ), .b(\ILAB0102.net17707 ), .c(\ILAB0102.net15728 ), .y(\ILAB0102.ILE1506.net2656 ));
  xci2_and3ftt _238_ ( .a(\ILAB0102.ILE1605.net0562 ), .b(\ILAB0102.net26482 ), .c(\net18572<1> ), .y(\ILAB0102.ILE1605.net2656 ));
  xci2_mux2h _239_ ( .a(\ILAB0102.net25628 ), .b(\ILAB0102.ILE1604.net0558 ), .s(\net18588<5> ), .y(\ILAB0102.ILE1604.net0541 ));
  xci2_ao21 _240_ ( .a(\net18584<2> ), .b(\ILAB0102.Clk_LAB<3> ), .c(\ILAB0102.net15889 ), .y(\ILAB0102.ILE1505.net2656 ));
  xci2_ao21 _241_ ( .a(\ILAB0102.net21128 ), .b(\ILAB0102.net25627 ), .c(\ILAB0102.net25061 ), .y(\ILAB0102.ILE1407.net2656 ));
  xci2_ao21ttf _242_ ( .a(\net18564<1> ), .b(\ILAB0202.net19732 ), .c(\ILAB0102.net16177 ), .y(\ILAB0102.ILE1508.net2656 ));
  xci2_ao21 _243_ ( .a(\net18532<1> ), .b(\ILAB0102.net22028 ), .c(\ILAB0102.net19642 ), .y(\ILAB0102.ILE1516.net2656 ));
  xci2_and3 _244_ ( .a(\ILAB0102.net17912 ), .b(\ILAB0102.net23243 ), .c(\net10391<0> ), .y(\ILAB0102.ILE1316.net2656 ));
  xci2_ao21 _245_ ( .a(\net10391<5> ), .b(\net10387<6> ), .c(\net10391<4> ), .y(\ILAB0103.ILE1301.net2656 ));
  xci2_and3 _246_ ( .a(\net10391<1> ), .b(\ILAB0102.net22207 ), .c(\net10391<0> ), .y(\ILAB0102.ILE1315.net2656 ));
  xci2_ao21 _247_ ( .a(\net10387<1> ), .b(\ILAB0102.net19372 ), .c(\net18536<0> ), .y(\ILAB0102.ILE1415.net2656 ));
  xci2_and3ftt _248_ ( .a(\ILAB0102.net16628 ), .b(\ILAB0102.net15754 ), .c(\ILAB0102.net25069 ), .y(\ILAB0102.ILE1305.net2656 ));
  xci2_mux2h _249_ ( .a(\ILAB0102.net20812 ), .b(\ILAB0102.ILE1604.net0558 ), .s(\net18588<1> ), .y(\ILAB0102.ILE1404.net2656 ));
  xci2_ao21 _250_ ( .a(\net18584<1> ), .b(\ILAB0102.net25629 ), .c(\ILAB0102.net25065 ), .y(\ILAB0102.ILE1405.net2656 ));
  xci2_ao21 _251_ ( .a(\ILAB0102.net23109 ), .b(\ILAB0102.net20029 ), .c(\ILAB0102.net15934 ), .y(\ILAB0102.ILE1005.net2656 ));
  xci2_and3fft _252_ ( .a(\ILAB0401.ILE0811.net01345 ), .b(\ILAB0401.Clk_LAB<3> ), .c(\ILAB0401.net23044 ), .y(\ILAB0401.ILE0811.net2656 ));
  xci2_nand3fft _253_ ( .a(\ILAB0401.net19914 ), .b(\ILAB0401.Clk_LAB<1> ), .c(\ILAB0401.net23494 ), .y(\ILAB0401.ILE0812.net2656 ));
  xci2_nor2 _254_ ( .a(\ILAB0401.net22657 ), .b(\ILAB0401.net16312 ), .y(\ILAB0401.ILE1012.net2656 ));
  xci2_nand3ftt _255_ ( .a(\ILAB0401.ILE0713.net0560 ), .b(\ILAB0401.net24143 ), .c(\ILAB0401.net21694 ), .y(\ILAB0401.ILE0712.net2656 ));
  xci2_and2ft _256_ ( .a(\ILAB0401.net22144 ), .b(\ILAB0401.net23784 ), .y(\ILAB0401.ILE0414.net2656 ));
  xci2_and2 _257_ ( .a(\ILAB0401.net19309 ), .b(\net16312<3> ), .y(\ILAB0401.ILE0516.net2656 ));
  xci2_nand3 _258_ ( .a(\ILAB0401.net22414 ), .b(\ILAB0401.net18904 ), .c(\ILAB0401.net19057 ), .y(\ILAB0401.ILE0514.net2656 ));
  xci2_nand2ft _259_ ( .a(\net16304<0> ), .b(\net16312<1> ), .y(\ILAB0401.ILE0515.net2656 ));
  xci2_ao21ftf _260_ ( .a(\net16271<6> ), .b(\ILAB0401.net19804 ), .c(\net11344<1> ), .y(\ILAB0401.ILE0115.net2656 ));
  xci2_and2 _261_ ( .a(\net11344<1> ), .b(\ILAB0401.ILE0116.net01339 ), .y(\ILAB0401.ILE0116.net2656 ));
  xci2_mux2h _262_ ( .a(\ILAB0401.net23197 ), .b(\ILAB0401.net21892 ), .s(\ILAB0401.net22254 ), .y(\ILAB0401.ILE0114.net2656 ));
  xci2_xnor2 _263_ ( .a(\ILAB0401.ILE0214.net01339 ), .b(\ILAB0401.net19939 ), .y(\ILAB0401.ILE0412.net2656 ));
  xci2_and3 _264_ ( .a(\ILAB0401.net18311 ), .b(\ILAB0401.net18315 ), .c(\ILAB0401.net19057 ), .y(\ILAB0401.ILE0513.net2656 ));
  xci2_and3 _264__1 ( .a(\ILAB0401.net18311 ), .b(\ILAB0401.net18315 ), .c(\ILAB0401.net19057 ), .y(\ILAB0401.ILE0513.net0541 ));
  xci2_nand3fft _265_ ( .a(\ILAB0401.net19350 ), .b(\ILAB0401.net18677 ), .c(\ILAB0401.net19174 ), .y(\ILAB0401.ILE0613.net2656 ));
  xci2_nand3fft _265__1 ( .a(\ILAB0401.net19350 ), .b(\ILAB0401.net18677 ), .c(\ILAB0401.net19174 ), .y(\ILAB0401.ILE0613.net0541 ));
  xci2_ao21 _266_ ( .a(\ILAB0401.net19174 ), .b(\ILAB0401.ILE0612.net01342 ), .c(\ILAB0401.net18949 ), .y(\ILAB0401.ILE0612.net2656 ));
  xci2_aoi21 _267_ ( .a(\ILAB0401.net23917 ), .b(\ILAB0401.net19714 ), .c(\ILAB0401.net18679 ), .y(\ILAB0401.ILE0512.net2656 ));
  xci2_ao21 _268_ ( .a(\net16283<3> ), .b(\ILAB0401.net21892 ), .c(\ILAB0401.net19084 ), .y(\ILAB0401.ILE0212.net2656 ));
  xci2_nand3ftt _269_ ( .a(\ILAB0401.net23648 ), .b(\ILAB0401.net24907 ), .c(\ILAB0401.ILE0214.net01339 ), .y(\ILAB0401.ILE0214.net2656 ));
  xci2_xnor2 _270_ ( .a(\ILAB0401.net23177 ), .b(\ILAB0401.net25537 ), .y(\ILAB0401.ILE0213.net2656 ));
  xci2_and3 _271_ ( .a(\net16304<5> ), .b(\ILAB0402.net20587 ), .c(\net16304<0> ), .y(\ILAB0402.ILE0701.net0541 ));
  xci2_and3 _272_ ( .a(\ILAB0401.net24549 ), .b(\ILAB0401.net24907 ), .c(\ILAB0401.net23153 ), .y(\ILAB0401.ILE0315.net2656 ));
  xci2_and3 _272__1 ( .a(\ILAB0401.net24549 ), .b(\ILAB0401.net24907 ), .c(\ILAB0401.net23153 ), .y(\ILAB0401.ILE0315.net0541 ));
  xci2_and3fft _273_ ( .a(\ILAB0401.net19309 ), .b(\ILAB0402.ILE0301.net01339 ), .c(\net16312<5> ), .y(\ILAB0402.ILE0301.net2656 ));
  xci2_nand2 _274_ ( .a(\ILAB0401.net22365 ), .b(\net16320<2> ), .y(\ILAB0401.ILE0415.net2656 ));
  xci2_nand3fft _275_ ( .a(\ILAB0401.net19174 ), .b(\ILAB0401.net18677 ), .c(\ILAB0401.net19238 ), .y(\ILAB0401.ILE0614.net2656 ));
  xci2_nand3fft _275__1 ( .a(\ILAB0401.net19174 ), .b(\ILAB0401.net18677 ), .c(\ILAB0401.net19238 ), .y(\ILAB0401.ILE0614.net0541 ));
  xci2_nand2 _276_ ( .a(\ILAB0401.net23964 ), .b(\ILAB0401.ILE0715.net01339 ), .y(\ILAB0401.ILE0715.net2656 ));
  xci2_nand3 _277_ ( .a(\ILAB0401.net22189 ), .b(\ILAB0401.net19328 ), .c(\ILAB0401.net22119 ), .y(\ILAB0401.ILE0615.net2656 ));
  xci2_and2 _278_ ( .a(\ILAB0401.net19309 ), .b(\net16320<3> ), .y(\ILAB0401.ILE0316.net2656 ));
  xci2_and2 _278__1 ( .a(\ILAB0401.net19309 ), .b(\net16320<3> ), .y(\ILAB0401.ILE0316.net0541 ));
  xci2_xnor2ft _279_ ( .a(\ILAB0401.net19309 ), .b(\ILAB0401.ILE0416.net01342 ), .y(\ILAB0401.ILE0416.net2656 ));
  xci2_ao21 _280_ ( .a(\net16308<2> ), .b(\ILAB0401.net17464 ), .c(\ILAB0401.ILE0616.net0558 ), .y(\ILAB0401.ILE0616.net2656 ));
  xci2_and3 _281_ ( .a(\net16312<5> ), .b(\net16312<0> ), .c(\net16304<0> ), .y(\ILAB0402.ILE0501.net2656 ));
  xci2_xnor2ft _282_ ( .a(\ILAB0402.ILE0401.net0558 ), .b(\ILAB0402.ILE0401.net01342 ), .y(\ILAB0402.ILE0401.net2656 ));
  xci2_ao21 _283_ ( .a(\net16308<3> ), .b(\ILAB0402.net20612 ), .c(\ILAB0402.net20929 ), .y(\ILAB0402.ILE0601.net0541 ));
  xci2_nand3ftt _284_ ( .a(\ILAB0401.net17014 ), .b(\net16267<3> ), .c(\net11247<1> ), .y(\ILAB0401.ILE0216.net2656 ));
  xci2_xnor2 _285_ ( .a(\net16324<1> ), .b(\net16324<4> ), .y(\ILAB0402.ILE0201.net2656 ));
  xci2_ao21 _286_ ( .a(\net16328<1> ), .b(\net11344<1> ), .c(\net11340<3> ), .y(\ILAB0402.ILE0101.net2656 ));
  xci2_nand3ftt _287_ ( .a(\ILAB0102.net26554 ), .b(\ILAB0102.net26329 ), .c(\ILAB0102.ILE1301.net01342 ), .y(\ILAB0102.ILE1302.net2656 ));
  xci2_mux2h _288_ ( .a(\net17198<6> ), .b(\net17202<4> ), .s(\ILAB0102.net26599 ), .y(\ILAB0102.ILE0901.net2656 ));
  xci2_and3fft _289_ ( .a(\ILAB0401.net23044 ), .b(\ILAB0401.net25312 ), .c(\ILAB0401.net18472 ), .y(\ILAB0401.ILE0911.net2656 ));
  xci2_and3fft _289__1 ( .a(\ILAB0401.net23044 ), .b(\ILAB0401.net25312 ), .c(\ILAB0401.net18472 ), .y(\ILAB0401.ILE0911.net0541 ));
  xci2_and2 _290_ ( .a(\ILAB0401.net21669 ), .b(\ILAB0401.net25494 ), .y(\ILAB0401.ILE1013.net2656 ));
  xci2_and3fft _291_ ( .a(\ILAB0401.net24979 ), .b(\ILAB0401.net24322 ), .c(\ILAB0401.ILE1010.net01342 ), .y(\ILAB0401.ILE1010.net2656 ));
  xci2_nand3fft _292_ ( .a(\ILAB0401.net18653 ), .b(\ILAB0401.net24885 ), .c(\ILAB0401.net21694 ), .y(\ILAB0401.ILE0912.net2656 ));
  xci2_and3fft _293_ ( .a(\ILAB0401.net21424 ), .b(\ILAB0401.net24977 ), .c(\ILAB0401.net18924 ), .y(\ILAB0401.ILE0913.net2656 ));
  xci2_nand3fft _294_ ( .a(\ILAB0401.net26078 ), .b(\ILAB0401.ILE0713.net0560 ), .c(\ILAB0401.net18992 ), .y(\ILAB0401.ILE0713.net2656 ));
  xci2_oa21 _295_ ( .a(\ILAB0401.net19913 ), .b(\ILAB0401.net22412 ), .c(\ILAB0401.ILE0714.net01339 ), .y(\ILAB0401.ILE0714.net0541 ));
  xci2_nand3 _296_ ( .a(\ILAB0401.net25519 ), .b(\ILAB0401.net21559 ), .c(\ILAB0401.ILE0813.net01339 ), .y(\ILAB0401.ILE0813.net2656 ));
  xci2_and3ftt _297_ ( .a(\ILAB0401.net24979 ), .b(\ILAB0401.net24322 ), .c(\ILAB0401.net22680 ), .y(\ILAB0401.ILE1011.net2656 ));
  xci2_nand3fft _298_ ( .a(\ILAB0401.net23042 ), .b(\ILAB0401.net22388 ), .c(\ILAB0401.net18922 ), .y(\ILAB0401.ILE0914.net2656 ));
  xci2_and3 _299_ ( .a(\ILAB0401.net24979 ), .b(\ILAB0401.Clk_LAB<2> ), .c(\ILAB0401.net25313 ), .y(\ILAB0401.ILE0910.net2656 ));
  xci2_nand3 _300_ ( .a(\ILAB0401.net19174 ), .b(\ILAB0401.net18499 ), .c(\ILAB0401.net20363 ), .y(\ILAB0401.ILE0611.net2656 ));
  xci2_aoi21 _301_ ( .a(\ILAB0401.net17977 ), .b(\ILAB0401.net24889 ), .c(\ILAB0401.net23719 ), .y(\ILAB0401.ILE0810.net0541 ));
  xci2_nand3 _302_ ( .a(\ILAB0401.net15637 ), .b(\ILAB0401.net21514 ), .c(\ILAB0401.ILE0711.net0558 ), .y(\ILAB0401.ILE0711.net2656 ));
  xci2_mux2h _303_ ( .a(\ILAB0201.net25897 ), .b(\ILAB0201.ILE0316.net01339 ), .s(\ILAB0201.net19354 ), .y(\ILAB0201.ILE0313.net2656 ));
  xci2_mux2h _304_ ( .a(\ILAB0102.net15709 ), .b(\ILAB0102.net17687 ), .s(\ILAB0102.net25114 ), .y(\ILAB0102.ILE0503.net2656 ));
  xci2_mux2h _305_ ( .a(\ILAB0102.net24142 ), .b(\ILAB0102.net19913 ), .s(\ILAB0102.net21488 ), .y(\ILAB0102.ILE0713.net2656 ));
  xci2_mux2h _306_ ( .a(\ILAB0102.net23494 ), .b(\ILAB0102.net22189 ), .s(\ILAB0102.net22099 ), .y(\ILAB0102.ILE0615.net2656 ));
  xci2_mux2h _307_ ( .a(\ILAB0103.net16556 ), .b(\ILAB0103.net26618 ), .s(\ILAB0103.net20452 ), .y(\ILAB0103.ILE1003.net2656 ));
  xci2_mux2h _308_ ( .a(\ILAB0103.net26194 ), .b(\ILAB0103.net26644 ), .s(\ILAB0102.net18922 ), .y(\ILAB0103.ILE0702.net2656 ));
  xci2_mux2h _309_ ( .a(\ILAB0103.net26149 ), .b(\ILAB0103.net20633 ), .s(\ILAB0103.net20522 ), .y(\ILAB0103.ILE0502.net2656 ));
  xci2_mux2h _310_ ( .a(\ILAB0102.net24527 ), .b(\ILAB0103.net26168 ), .s(\ILAB0103.net20299 ), .y(\ILAB0103.ILE0903.net2656 ));
  xci2_mux2h _311_ ( .a(\ILAB0103.net26192 ), .b(\ILAB0103.net26438 ), .s(\ILAB0103.net20299 ), .y(\ILAB0103.ILE0703.net2656 ));
  xci2_mux2h _312_ ( .a(\ILAB0102.net24212 ), .b(\ILAB0103.net20612 ), .s(\ILAB0103.net20614 ), .y(\ILAB0103.ILE0501.net2656 ));
  xci2_mux2h _313_ ( .a(\ILAB0102.ILE0711.net0562 ), .b(\ILAB0102.net22684 ), .s(\ILAB0102.net25159 ), .y(\ILAB0102.ILE0711.net2656 ));
  xci2_mux2h _314_ ( .a(\ILAB0102.net25609 ), .b(\ILAB0102.net25020 ), .s(\ILAB0102.net25114 ), .y(\ILAB0102.ILE0504.net2656 ));
  xci2_mux2h _315_ ( .a(\ILAB0102.net26689 ), .b(\ILAB0102.net20678 ), .s(\ILAB0102.net25114 ), .y(\ILAB0102.ILE0802.net2656 ));
  xci2_mux2h _316_ ( .a(\ILAB0102.net26149 ), .b(\ILAB0102.net20588 ), .s(\ILAB0102.net25114 ), .y(\ILAB0102.ILE0602.net2656 ));
  xci2_mux2h _317_ ( .a(\ILAB0102.ILE0604.net0562 ), .b(\ILAB0102.net17663 ), .s(\ILAB0102.net25114 ), .y(\ILAB0102.ILE0604.net2656 ));
  xci2_mux2h _318_ ( .a(\ILAB0102.net15817 ), .b(\ILAB0102.net18229 ), .s(\ILAB0102.net18634 ), .y(\ILAB0102.ILE0706.net2656 ));
  xci2_mux2h _319_ ( .a(\ILAB0102.net21062 ), .b(\ILAB0102.net19620 ), .s(\ILAB0102.net19624 ), .y(\ILAB0102.ILE0608.net2656 ));
  xci2_mux2h _320_ ( .a(\ILAB0102.net24889 ), .b(\ILAB0102.net24165 ), .s(\ILAB0102.net25159 ), .y(\ILAB0102.ILE0710.net2656 ));
  xci2_mux2h _321_ ( .a(\ILAB0102.net24752 ), .b(\ILAB0102.net24863 ), .s(\ILAB0102.net16222 ), .y(\ILAB0102.ILE1011.net2656 ));
  xci2_mux2h _322_ ( .a(\ILAB0102.net21152 ), .b(\ILAB0102.net15908 ), .s(\ILAB0102.net25133 ), .y(\ILAB0102.ILE1306.net2656 ));
  xci2_mux2h _323_ ( .a(\net18564<1> ), .b(\net10337<3> ), .s(\ILAB0102.net16222 ), .y(\ILAB0102.ILE1312.net2656 ));
  xci2_mux2h _324_ ( .a(\ILAB0103.net26574 ), .b(\ILAB0103.net26573 ), .s(\ILAB0103.net20452 ), .y(\ILAB0103.ILE1203.net2656 ));
  xci2_mux2h _325_ ( .a(\ILAB0103.net26329 ), .b(\ILAB0103.net16583 ), .s(\net10399<5> ), .y(\ILAB0103.ILE1102.net2656 ));
  xci2_mux2h _326_ ( .a(\ILAB0102.net19847 ), .b(\ILAB0102.net21352 ), .s(\net10391<0> ), .y(\ILAB0102.ILE1215.net2656 ));
  xci2_mux2h _327_ ( .a(\ILAB0102.net17977 ), .b(\ILAB0102.net17617 ), .s(\ILAB0102.net18679 ), .y(\ILAB0102.ILE0812.net2656 ));
  xci2_mux2h _328_ ( .a(\net16275<6> ), .b(\net11344<3> ), .s(\ILAB0302.net20569 ), .y(\ILAB0302.ILE1601.net2656 ));
  xci2_xnor2 _329_ ( .a(\Fast_out_28<0> ), .b(\ILAB0102.net21064 ), .y(\ILAB0102.ILE0408.net2656 ));
  xci2_xnor2 _330_ ( .a(\ILAB0102.net17509 ), .b(\ILAB0102.net19309 ), .y(\ILAB0102.ILE0616.net2656 ));
  xci2_xnor2 _331_ ( .a(\ILAB0102.ILE0416.net0558 ), .b(\ILAB0102.net17014 ), .y(\ILAB0102.ILE0416.net2656 ));
  xci2_xnor2 _332_ ( .a(\net10430<6> ), .b(\ILAB0102.net26754 ), .y(\ILAB0102.ILE0203.net2656 ));
  xci2_xnor2 _333_ ( .a(\ILAB0102.net18589 ), .b(\Fast_out_28<2> ), .y(\ILAB0102.ILE0506.net2656 ));
  xci2_xnor2 _334_ ( .a(\ILAB0102.net15799 ), .b(\ILAB0102.net15844 ), .y(\ILAB0102.ILE0405.net2656 ));
  xci2_xnor2 _335_ ( .a(\ILAB0103.ILE0402.net0558 ), .b(\net10427<3> ), .y(\ILAB0103.ILE0402.net2656 ));
  xci2_xnor2 _336_ ( .a(\ILAB0103.net25114 ), .b(\ILAB0103.net25989 ), .y(\ILAB0103.ILE0605.net2656 ));
  xci2_xnor2 _337_ ( .a(\ILAB0102.net20612 ), .b(\ILAB0102.net20724 ), .y(\ILAB0102.ILE0402.net2656 ));
  xci2_xnor2 _338_ ( .a(\ILAB0102.net20929 ), .b(\ILAB0102.net20634 ), .y(\ILAB0102.ILE0502.net2656 ));
  xci2_xnor2 _339_ ( .a(\net10426<6> ), .b(\ILAB0102.net26014 ), .y(\ILAB0102.ILE0304.net2656 ));
  xci2_xnor2 _340_ ( .a(\net11487<6> ), .b(\net10431<3> ), .y(\ILAB0103.ILE0302.net2656 ));
  xci2_xnor2 _341_ ( .a(\ILAB0102.net22549 ), .b(\ILAB0102.net19804 ), .y(\ILAB0102.ILE0414.net2656 ));
  xci2_xnor2 _342_ ( .a(\ILAB0102.net24124 ), .b(\ILAB0102.net23895 ), .y(\ILAB0102.ILE0410.net2656 ));
  xci2_and2 _343_ ( .a(\ILAB0102.net23872 ), .b(\ILAB0102.net23874 ), .y(\ILAB0102.ILE0411.net2656 ));
  xci2_and3 _344_ ( .a(\ILAB0102.net17753 ), .b(\ILAB0102.net20182 ), .c(\ILAB0102.net18112 ), .y(\ILAB0102.ILE0407.net2656 ));
  xci2_xnor2 _345_ ( .a(\ILAB0103.net16114 ), .b(\Fast_out_29<4> ), .y(\ILAB0103.ILE0504.net2656 ));
  xci2_xnor2 _346_ ( .a(\ILAB0103.net23132 ), .b(\ILAB0103.net25584 ), .y(\ILAB0103.ILE0805.net2656 ));
  xci2_xnor2 _347_ ( .a(\ILAB0102.net21694 ), .b(\ILAB0102.net19935 ), .y(\ILAB0102.ILE0712.net2656 ));
  xci2_and2 _348_ ( .a(\ILAB0103.net17374 ), .b(\ILAB0103.net20497 ), .y(\ILAB0103.ILE0705.net2656 ));
  xci2_and3 _349_ ( .a(\ILAB0103.net15799 ), .b(\ILAB0103.net24999 ), .c(\ILAB0103.net15844 ), .y(\ILAB0103.ILE0505.net2656 ));
  xci2_xnor2 _350_ ( .a(\ILAB0102.ILE0510.net0558 ), .b(\ILAB0102.net16762 ), .y(\ILAB0102.ILE0510.net2656 ));
  xci2_xnor2 _351_ ( .a(\ILAB0102.net25969 ), .b(\ILAB0102.net25249 ), .y(\ILAB0102.ILE0607.net2656 ));
  xci2_and3 _352_ ( .a(\ILAB0102.net18744 ), .b(\ILAB0102.net25448 ), .c(\ILAB0102.net17102 ), .y(\ILAB0102.ILE0507.net2656 ));
  xci2_and2 _353_ ( .a(\ILAB0102.net19463 ), .b(\ILAB0102.net16763 ), .y(\ILAB0102.ILE0509.net2656 ));
  xci2_and3 _354_ ( .a(\ILAB0102.net16672 ), .b(\ILAB0102.net25447 ), .c(\ILAB0102.net19129 ), .y(\ILAB0102.ILE0409.net2656 ));
  xci2_xnor2 _355_ ( .a(\ILAB0102.net19939 ), .b(\ILAB0102.net23175 ), .y(\ILAB0102.ILE0313.net2656 ));
  xci2_and2 _356_ ( .a(\ILAB0102.net19013 ), .b(\ILAB0102.net26100 ), .y(\ILAB0102.ILE0413.net2656 ));
  xci2_and3 _357_ ( .a(\ILAB0102.net19417 ), .b(\ILAB0102.net19867 ), .c(\ILAB0102.net19868 ), .y(\ILAB0102.ILE0412.net2656 ));
  xci2_xnor2 _358_ ( .a(\net11487<3> ), .b(\ELLR15_28<3> ), .y(\ILAB0102.ILE0216.net2656 ));
  xci2_and2 _359_ ( .a(\ILAB0102.net23287 ), .b(\ILAB0102.net22297 ), .y(\ILAB0102.ILE0215.net2656 ));
  xci2_xnor2 _360_ ( .a(\net11495<6> ), .b(\ILAB0103.net17865 ), .y(\ILAB0103.ILE0301.net2656 ));
  xci2_and3 _361_ ( .a(\net10431<1> ), .b(\ELLR14_28<3> ), .c(\net10431<0> ), .y(\ILAB0102.ILE0315.net2656 ));
  xci2_xnor2 _362_ ( .a(\ILAB0102.ILE0613.net0558 ), .b(\ILAB0102.net25519 ), .y(\ILAB0102.ILE0613.net2656 ));
  xci2_xnor2 _363_ ( .a(\net10419<5> ), .b(\ILAB0103.net20524 ), .y(\ILAB0103.ILE0601.net2656 ));
  xci2_and3 _364_ ( .a(\ILAB0102.net19687 ), .b(\ILAB0102.net19329 ), .c(\net10419<0> ), .y(\ILAB0102.ILE0614.net2656 ));
  xci2_and2 _365_ ( .a(\ILAB0102.net15367 ), .b(\ILAB0102.net22144 ), .y(\ILAB0102.ILE0311.net2656 ));
  xci2_and3 _366_ ( .a(\ILAB0102.net19084 ), .b(\ILAB0102.net23377 ), .c(\ILAB0102.net23379 ), .y(\ILAB0102.ILE0312.net2656 ));
  xci2_nand2 _367_ ( .a(\ILAB0102.net18407 ), .b(\ILAB0102.net25852 ), .y(\ILAB0102.ILE0309.net2656 ));
  xci2_dffcl _368_ ( .d(\ILAB0102.net26509 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE1501.net01339 ), .q(\ILAB0102.ILE1502.net2656 ));
  xci2_dffcl _369_ ( .d(\ILAB0102.net24664 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net26124 ), .q(\ILAB0102.ILE0806.net2656 ));
  xci2_dffcl _370_ ( .d(\ILAB0102.net23269 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE1216.net01339 ), .q(\ILAB0102.ILE1014.net2656 ));
  xci2_dffcl _370__1 ( .d(\ILAB0102.net23269 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE1216.net01339 ), .q(\ILAB0102.ILE1014.net0541 ));
  xci2_dffcl _371_ ( .d(\ILAB0102.net21197 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.Clk_LAB<1> ), .q(\ILAB0103.ILE1002.net0541 ));
  xci2_dffcl _372_ ( .d(\ILAB0103.net15504 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.net15502 ), .q(\ILAB0103.ILE1202.net2656 ));
  xci2_dffcl _373_ ( .d(\ILAB0103.net20679 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0102.ILE1216.net01339 ), .q(\ILAB0103.ILE0802.net2656 ));
  xci2_dffcl _374_ ( .d(\ILAB0102.net21667 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE1416.net01339 ), .q(\ILAB0102.ILE1015.net2656 ));
  xci2_dffcl _375_ ( .d(\net10407<6> ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.Clk_LAB<1> ), .q(\ILAB0103.ILE0902.net2656 ));
  xci2_dffcl _376_ ( .d(\ILAB0102.net22097 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0716.net01339 ), .q(\ILAB0102.ILE0715.net2656 ));
  xci2_dffcl _376__1 ( .d(\ILAB0102.net22097 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0716.net01339 ), .q(\ILAB0102.ILE0715.net0541 ));
  xci2_dffcl _377_ ( .d(\ILAB0102.net17618 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0516.net01339 ), .q(\ILAB0102.ILE0810.net2656 ));
  xci2_dffcl _377__1 ( .d(\ILAB0102.net17618 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0516.net01339 ), .q(\ILAB0102.ILE0810.net0541 ));
  xci2_dffcl _378_ ( .d(\ILAB0102.net25830 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net17194 ), .q(\ILAB0102.ILE1007.net2656 ));
  xci2_dffcl _379_ ( .d(\net17194<3> ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE1101.net01339 ), .q(\ILAB0102.ILE1102.net2656 ));
  xci2_dffcl _379__1 ( .d(\net17194<3> ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE1101.net01339 ), .q(\ILAB0102.ILE1102.net0541 ));
  xci2_dffcl _380_ ( .d(\net17202<3> ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net26124 ), .q(\ILAB0102.ILE0902.net2656 ));
  xci2_dffcl _381_ ( .d(\ILAB0102.net20344 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE1001.net01345 ), .q(\ILAB0102.ILE0703.net2656 ));
  xci2_dffcl _381__1 ( .d(\ILAB0102.net20344 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE1001.net01345 ), .q(\ILAB0102.ILE0703.net0541 ));
  xci2_dffcl _382_ ( .d(\ILAB0102.net17374 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE1001.net01345 ), .q(\ILAB0102.ILE0705.net2656 ));
  xci2_dffcl _383_ ( .d(\ILAB0102.net18002 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net19462 ), .q(\ILAB0102.ILE0708.net2656 ));
  xci2_dffcl _384_ ( .d(\ILAB0102.net25314 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0516.net01339 ), .q(\ILAB0102.ILE0910.net2656 ));
  xci2_dffcl _385_ ( .d(\ILAB0102.net24079 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net16267 ), .q(\ILAB0102.ILE1210.net2656 ));
  xci2_dffcl _386_ ( .d(\ILAB0102.net18184 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0202.ILE0106.net01339 ), .q(\ILAB0102.ILE1406.net2656 ));
  xci2_dffcl _387_ ( .d(\ILAB0102.net25764 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0202.ILE0108.net01339 ), .q(\ILAB0102.ILE1408.net2656 ));
  xci2_dffcl _388_ ( .d(\ILAB0102.net18814 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE1416.net01339 ), .q(\ILAB0102.ILE1416.net2656 ));
  xci2_dffcl _389_ ( .d(\ILAB0103.net20454 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.ILE1602.net0560 ), .q(\ILAB0103.ILE1302.net2656 ));
  xci2_dffcl _390_ ( .d(\ILAB0102.net20407 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE1416.net01339 ), .q(\ILAB0102.ILE1414.net2656 ));
  xci2_dffcl _391_ ( .d(\ILAB0102.net16537 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net25988 ), .q(\ILAB0102.ILE1004.net2656 ));
  xci2_dffcl _392_ ( .d(\ILAB0401.net25267 ), .clk(\ILAB0401.Clk_LAB<0> ), .clr(\ILAB0401.ILE0113.net01339 ), .q(\ILAB0401.ILE0113.net2656 ));
  xci2_dffcl _392__1 ( .d(\ILAB0401.net25267 ), .clk(\ILAB0401.Clk_LAB<0> ), .clr(\ILAB0401.ILE0113.net01339 ), .q(\ILAB0401.ILE0113.net0541 ));
  xci2_dffcl _393_ ( .d(\ILAB0401.net24930 ), .clk(\ILAB0401.Clk_LAB<0> ), .clr(\ILAB0401.net23377 ), .q(\ILAB0401.ILE0312.net2656 ));
  xci2_dffcl _393__1 ( .d(\ILAB0401.net24930 ), .clk(\ILAB0401.Clk_LAB<0> ), .clr(\ILAB0401.net23377 ), .q(\ILAB0401.ILE0312.net0541 ));
  xci2_dffcl _394_ ( .d(\ILAB0401.net23175 ), .clk(\ILAB0401.Clk_LAB<0> ), .clr(\net16279<6> ), .q(\ILAB0401.ILE0313.net2656 ));
  xci2_dffcl _395_ ( .d(\ILAB0401.net21604 ), .clk(\ILAB0401.Clk_LAB<0> ), .clr(\ILAB0401.ILE0716.net01339 ), .q(\ILAB0401.ILE0716.net2656 ));
  xci2_dffcl _396_ ( .d(\ILAB0402.ILE0502.net0562 ), .clk(\ILAB0402.Clk_LAB<1> ), .clr(\ILAB0401.ILE0716.net01339 ), .q(\ILAB0402.ILE0502.net2656 ));
  xci2_dffcl _396__1 ( .d(\ILAB0402.ILE0502.net0562 ), .clk(\ILAB0402.Clk_LAB<1> ), .clr(\ILAB0401.ILE0716.net01339 ), .q(\ILAB0402.ILE0502.net0541 ));
  xci2_dffcl _397_ ( .d(\ILAB0402.net16944 ), .clk(\ILAB0402.Clk_LAB<1> ), .clr(\ILAB0402.net26775 ), .q(\ILAB0402.ILE0202.net2656 ));
  xci2_dffcl _397__1 ( .d(\ILAB0402.net16944 ), .clk(\ILAB0402.Clk_LAB<1> ), .clr(\ILAB0402.net26775 ), .q(\ILAB0402.ILE0202.net0541 ));
  xci2_dffcl _398_ ( .d(\ILAB0402.net16719 ), .clk(\ILAB0402.Clk_LAB<1> ), .clr(\ILAB0402.ILE0102.net01339 ), .q(\ILAB0402.ILE0102.net2656 ));
  xci2_dffcl _398__1 ( .d(\ILAB0402.net16719 ), .clk(\ILAB0402.Clk_LAB<1> ), .clr(\ILAB0402.ILE0102.net01339 ), .q(\ILAB0402.ILE0102.net0541 ));
  xci2_dff _399_ ( .d(\net17202<0> ), .clk(\ILAB0101.Clk_LAB<0> ), .q(\ILAB0101.ILE0916.net2656 ));
  xci2_dff _399__1 ( .d(\net17202<0> ), .clk(\ILAB0101.Clk_LAB<0> ), .q(\ILAB0101.ILE0916.net0541 ));
  xci2_dffcl _400_ ( .d(\ILAB0401.net22524 ), .clk(\ILAB0401.Clk_LAB<0> ), .clr(\ILAB0401.ILE0816.net01342 ), .q(\ILAB0401.ILE0814.net2656 ));
  xci2_dffcl _400__1 ( .d(\ILAB0401.net22524 ), .clk(\ILAB0401.Clk_LAB<0> ), .clr(\ILAB0401.ILE0816.net01342 ), .q(\ILAB0401.ILE0814.net0541 ));
  xci2_dffcl _401_ ( .d(\ILAB0401.net23269 ), .clk(\ILAB0401.Clk_LAB<0> ), .clr(\ILAB0401.ILE0916.net01339 ), .q(\ILAB0401.ILE1014.net2656 ));
  xci2_dffcl _402_ ( .d(\ILAB0401.net17212 ), .clk(\ILAB0401.Clk_LAB<0> ), .clr(\ILAB0401.net21037 ), .q(\ILAB0401.ILE0710.net2656 ));
  xci2_dffcl _402__1 ( .d(\ILAB0401.net17212 ), .clk(\ILAB0401.Clk_LAB<0> ), .clr(\ILAB0401.net21037 ), .q(\ILAB0401.ILE0710.net0541 ));
  xci2_dffcl _403_ ( .d(\ILAB0201.net23154 ), .clk(\ILAB0201.Clk_LAB<0> ), .clr(\ILAB0201.ILE0316.net01345 ), .q(\ILAB0201.ILE0314.net2656 ));
  xci2_dffcl _404_ ( .d(\Fast_out_28<5> ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net20722 ), .q(\ILAB0102.ILE0403.net2656 ));
  xci2_dffcl _405_ ( .d(\ILAB0102.net19959 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0316.net01339 ), .q(\ILAB0102.ILE0714.net2656 ));
  xci2_dffcl _405__1 ( .d(\ILAB0102.net19959 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0316.net01339 ), .q(\ILAB0102.ILE0714.net0541 ));
  xci2_dffcl _406_ ( .d(\ILAB0102.net23989 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0516.net01339 ), .q(\ILAB0102.ILE0515.net2656 ));
  xci2_dffcl _406__1 ( .d(\ILAB0102.net23989 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0516.net01339 ), .q(\ILAB0102.ILE0515.net0541 ));
  xci2_dffcl _407_ ( .d(\ILAB0103.net17394 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.net15502 ), .q(\ILAB0103.ILE1004.net2656 ));
  xci2_dffcl _408_ ( .d(\ILAB0103.net26464 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.net26752 ), .q(\ILAB0103.ILE0602.net2656 ));
  xci2_dffcl _408__1 ( .d(\ILAB0103.net26464 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.net26752 ), .q(\ILAB0103.ILE0602.net0541 ));
  xci2_dffcl _409_ ( .d(\ILAB0103.net26259 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\net10423<6> ), .q(\ILAB0103.ILE0503.net2656 ));
  xci2_dffcl _409__1 ( .d(\ILAB0103.net26259 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\net10423<6> ), .q(\ILAB0103.ILE0503.net0541 ));
  xci2_dffcl _410_ ( .d(\ILAB0103.net20274 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.net15502 ), .q(\ILAB0103.ILE0904.net2656 ));
  xci2_dffcl _411_ ( .d(\ILAB0103.net15684 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.net26437 ), .q(\ILAB0103.ILE0704.net2656 ));
  xci2_dffcl _412_ ( .d(\Fast_out_29<7> ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.ILE0401.net01339 ), .q(\ILAB0103.ILE0401.net2656 ));
  xci2_dffcl _412__1 ( .d(\Fast_out_29<7> ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.ILE0401.net01339 ), .q(\ILAB0103.ILE0401.net0541 ));
  xci2_dffcl _413_ ( .d(\ILAB0102.net21514 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net19462 ), .q(\ILAB0102.ILE0611.net2656 ));
  xci2_dffcl _413__1 ( .d(\ILAB0102.net21514 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net19462 ), .q(\ILAB0102.ILE0611.net0541 ));
  xci2_dffcl _414_ ( .d(\Fast_out_28<4> ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net20722 ), .q(\ILAB0102.ILE0404.net2656 ));
  xci2_dffcl _415_ ( .d(\net17206<1> ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0801.net01339 ), .q(\ILAB0102.ILE0801.net2656 ));
  xci2_dffcl _415__1 ( .d(\net17206<1> ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0801.net01339 ), .q(\ILAB0102.ILE0801.net0541 ));
  xci2_dffcl _416_ ( .d(\net17214<5> ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0601.net01339 ), .q(\ILAB0102.ILE0601.net2656 ));
  xci2_dffcl _416__1 ( .d(\net17214<5> ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0601.net01339 ), .q(\ILAB0102.ILE0601.net0541 ));
  xci2_dffcl _417_ ( .d(\ILAB0102.net25989 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0801.net01339 ), .q(\ILAB0102.ILE0605.net2656 ));
  xci2_dffcl _418_ ( .d(\ILAB0102.net16069 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net26392 ), .q(\ILAB0102.ILE0606.net2656 ));
  xci2_dffcl _419_ ( .d(\ILAB0102.net19622 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net18004 ), .q(\ILAB0102.ILE0508.net2656 ));
  xci2_dffcl _420_ ( .d(\ILAB0102.net24169 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net18562 ), .q(\ILAB0102.ILE0610.net2656 ));
  xci2_dffcl _421_ ( .d(\ILAB0102.net22659 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net21690 ), .q(\ILAB0102.ILE1012.net2656 ));
  xci2_dffcl _422_ ( .d(\ILAB0102.net18699 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net25744 ), .q(\ILAB0102.ILE1307.net2656 ));
  xci2_dffcl _423_ ( .d(\ILAB0102.net21244 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net16267 ), .q(\ILAB0102.ILE1212.net2656 ));
  xci2_dffcl _424_ ( .d(\ILAB0103.net15594 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.net15502 ), .q(\ILAB0103.ILE1204.net2656 ));
  xci2_dffcl _425_ ( .d(\ILAB0103.net26664 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.Clk_LAB<1> ), .q(\ILAB0103.ILE1103.net2656 ));
  xci2_dffcl _426_ ( .d(\ILAB0102.net24414 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE1216.net01339 ), .q(\ILAB0102.ILE1216.net2656 ));
  xci2_dffcl _426__1 ( .d(\ILAB0102.net24414 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE1216.net01339 ), .q(\ILAB0102.ILE1216.net0541 ));
  xci2_dffcl _427_ ( .d(\ILAB0102.net18654 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net21559 ), .q(\ILAB0102.ILE0813.net2656 ));
  xci2_dffcl _428_ ( .d(\net11344<0> ), .clk(\ILAB0302.Clk_LAB<1> ), .clr(\ILAB0302.ILE1501.net01339 ), .q(\ILAB0302.ILE1501.net2656 ));
  xci2_dffcl _428__1 ( .d(\net11344<0> ), .clk(\ILAB0302.Clk_LAB<1> ), .clr(\ILAB0302.ILE1501.net01339 ), .q(\ILAB0302.ILE1501.net0541 ));
  xci2_dffcl _429_ ( .d(\ILAB1001.net25762 ), .clk(\ILAB1001.Clk_LAB<2> ), .clr(\ILAB1001.ILE1610.net0562 ), .q(\ILAB1001.ILE1410.net2656 ));
  xci2_dffcl _430_ ( .d(\net17226<1> ), .clk(\ILAB0101.Clk_LAB<0> ), .clr(\ILAB0101.ILE0216.net01339 ), .q(\ILAB0101.ILE0215.net0541 ));
  xci2_dffcl _431_ ( .d(\net10430<6> ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\net17230<6> ), .q(\ILAB0102.ILE0202.net2656 ));
  xci2_dffcl _432_ ( .d(\ILAB0102.net19913 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0516.net01339 ), .q(\ILAB0102.ILE0513.net2656 ));
  xci2_dffcl _433_ ( .d(\net10423<3> ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0516.net01339 ), .q(\ILAB0102.ILE0516.net2656 ));
  xci2_dffcl _434_ ( .d(\ILAB0103.net23134 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0102.ILE1216.net01339 ), .q(\ILAB0103.ILE0804.net2656 ));
  xci2_dffcl _435_ ( .d(\ILAB0103.ILE0701.net01345 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.ILE0701.net01339 ), .q(\ILAB0103.ILE0701.net2656 ));
  xci2_dffcl _436_ ( .d(\ILAB0103.net20162 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.net26214 ), .q(\ILAB0103.ILE0403.net2656 ));
  xci2_dffcl _437_ ( .d(\ILAB0103.net25114 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.net24997 ), .q(\ILAB0103.ILE0604.net2656 ));
  xci2_dffcl _438_ ( .d(\ILAB0103.net16114 ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.net20655 ), .q(\ILAB0103.ILE0404.net2656 ));
  xci2_dffcl _439_ ( .d(\net11495<6> ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0103.ILE0201.net01339 ), .q(\ILAB0103.ILE0201.net2656 ));
  xci2_dffcl _440_ ( .d(\ILAB0102.net21467 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net19462 ), .q(\ILAB0102.ILE0511.net2656 ));
  xci2_dffcl _441_ ( .d(\net10426<6> ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\net17230<6> ), .q(\ILAB0102.ILE0204.net2656 ));
  xci2_dffcl _442_ ( .d(\ILAB0102.net20704 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0501.net01339 ), .q(\ILAB0102.ILE0501.net2656 ));
  xci2_dffcl _443_ ( .d(\ILAB0102.net20614 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0401.net01339 ), .q(\ILAB0102.ILE0401.net2656 ));
  xci2_dffcl _444_ ( .d(\ILAB0102.net15799 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0601.net01339 ), .q(\ILAB0102.ILE0305.net2656 ));
  xci2_dffcl _445_ ( .d(\ILAB0102.net18589 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net15548 ), .q(\ILAB0102.ILE0406.net2656 ));
  xci2_dffcl _446_ ( .d(\Fast_out_28<0> ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net23332 ), .q(\ILAB0102.ILE0308.net2656 ));
  xci2_dffcl _447_ ( .d(\ILAB0102.net24124 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net25537 ), .q(\ILAB0102.ILE0310.net2656 ));
  xci2_dffcl _448_ ( .d(\ILAB0102.net18949 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0516.net01339 ), .q(\ILAB0102.ILE0612.net2656 ));
  xci2_dffcl _449_ ( .d(\ILAB0102.net25969 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net19462 ), .q(\ILAB0102.ILE0707.net2656 ));
  xci2_dffcl _450_ ( .d(\ILAB0102.net19939 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.net25537 ), .q(\ILAB0102.ILE0213.net2656 ));
  xci2_dffcl _451_ ( .d(\net11487<6> ), .clk(\ILAB0103.Clk_LAB<3> ), .clr(\ILAB0102.ILE0516.net01339 ), .q(\ILAB0103.ILE0303.net2656 ));
  xci2_dffcl _452_ ( .d(\net11487<3> ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0316.net01339 ), .q(\ILAB0102.ILE0316.net2656 ));
  xci2_dffcl _453_ ( .d(\ILAB0102.net17509 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0716.net01339 ), .q(\ILAB0102.ILE0716.net2656 ));
  xci2_dffcl _454_ ( .d(\ILAB0102.net17617 ), .clk(\ILAB0102.Clk_LAB<0> ), .clr(\ILAB0102.ILE0516.net01339 ), .q(\ILAB0102.ILE0514.net2656 ));
  mux2i_P_UCCLAB \IIO33.I0.I25  ( .d0(\IIO33.I0.net209 ), .d1(GND), .sl0(GND), .x(\IIO33.I0.net0153 ));
  invtd52_AVDD \IIO33.I0.I26  ( .a(\IIO33.I0.net0153 ), .en(VDD), .x(\LongBus_21<15> ));
  buftd52C_UCCLAB \I1803.I29  ( .a(\LongBus_21<15> ), .en(VDD), .x(\net8320<0> ));
  inv_4_UCCLAB \ILAB0401.ILE0916.I714  ( .a(\net8320<0> ), .x(\ILAB0401.ILE0916.net01345 ));
  mux2i_P_UCCLAB \IIO33.I0.I27  ( .d0(\IIO33.I0.net209 ), .d1(GND), .sl0(GND), .x(\IIO33.I0.net0151 ));
  invtd52_AVDD \IIO33.I0.I8  ( .a(\IIO33.I0.net0151 ), .en(VDD), .x(\LongBus_20<7> ));
  buftd52C_UCCLAB \I1804.I37  ( .a(\LongBus_20<7> ), .en(VDD), .x(\net8311<8> ));
  inv_4_UCCLAB \ILAB0401.ILE1601.I714  ( .a(\net8311<8> ), .x(\ILAB0401.ILE1601.net01345 ));
  inv_4_UCCLAB \ILAB0401.ILE1016.I713  ( .a(\net8320<0> ), .x(\ILAB0401.ILE1016.net01342 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0913.Ihi7  ( .en(GND), .in(\ILAB0401.ILE0916.net01345 ), .out(\ILAB0401.net25312 ));
  inv_8_UCCLAB \ILAB0401.ILE1601.I666  ( .a(\ILAB0401.ILE1601.net01345 ), .x(\net21156<0> ));
  buftd4_UCCLAB \ILAB0401.I236  ( .a(\net21156<0> ), .en(VDD), .x(\ILAB0401.net027166 ));
  mux2p_2_UCCLAB \ILAB0401.I5605.I4  ( .d0(\ILAB0401.net027166 ), .d1(GND), .s0(GND), .x(\ILAB0401.I5605.net25 ));
  invd16_seth_UCCLAB \ILAB0401.I5605.I5  ( .a(\ILAB0401.I5605.net25 ), .c(VDD), .x(\ILAB0401.Clk_int<1> ));
  mux2d1i_1_P_UCCLAB \ILAB0401.I5366.I79  ( .d0(\ILAB0401.Clk_int<1> ), .d1i(GND), .sl0(GND), .x(\ILAB0401.I5366.net0110 ));
  invd52_UCCLAB \ILAB0401.I5366.I75  ( .a(\ILAB0401.I5366.net0110 ), .x(\ILAB0401.net15299<2> ));
  invd32_UCCLAB \ILAB0401.I5591.I2  ( .a(\ILAB0401.net15299<2> ), .x(\ILAB0401.Clk_LAB<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE1013.Ihi7  ( .en(GND), .in(\ILAB0401.ILE1016.net01342 ), .out(\ILAB0401.net16312 ));
  buftd4_UCCLAB \ILAB0401.I238  ( .a(\net21156<0> ), .en(VDD), .x(\ILAB0401.net27188 ));
  mux2p_2_UCCLAB \ILAB0401.I5605.I0  ( .d0(\ILAB0401.net27188 ), .d1(GND), .s0(GND), .x(\ILAB0401.I5605.net29 ));
  invd16_seth_UCCLAB \ILAB0401.I5605.I1  ( .a(\ILAB0401.I5605.net29 ), .c(VDD), .x(\ILAB0401.Clk_int<3> ));
  mux2d1i_1_P_UCCLAB \ILAB0401.I5366.I81  ( .d0(\ILAB0401.Clk_int<3> ), .d1i(GND), .sl0(GND), .x(\ILAB0401.I5366.net0102 ));
  invd52_UCCLAB \ILAB0401.I5366.I77  ( .a(\ILAB0401.I5366.net0102 ), .x(\ILAB0401.net15299<0> ));
  invd32_UCCLAB \ILAB0401.I5591.I0  ( .a(\ILAB0401.net15299<0> ), .x(\ILAB0401.Clk_LAB<3> ));
  mux2i_P_UCCLAB \IIO33.I1.I25  ( .d0(\IIO33.I1.net209 ), .d1(GND), .sl0(GND), .x(\IIO33.I1.net0153 ));
  invtd52_AVDD \IIO33.I1.I26  ( .a(\IIO33.I1.net0153 ), .en(VDD), .x(\LongBus_21<14> ));
  buftd52C_UCCLAB \I1803.I26  ( .a(\LongBus_21<14> ), .en(VDD), .x(\net8320<1> ));
  buftd52C_UCCLAB \I3740.I26  ( .a(\net8320<1> ), .en(VDD), .x(\LongBus_78<14> ));
  inv_4_UCCLAB \ILAB0101.ILE1516.I714  ( .a(\LongBus_78<14> ), .x(\ILAB0101.ILE1516.net01345 ));
  mux2i_P_UCCLAB \IIO33.I2.I27  ( .d0(\IIO33.I2.net209 ), .d1(GND), .sl0(GND), .x(\IIO33.I2.net0151 ));
  mux2i_P_UCCLAB \IIO33.I2.I25  ( .d0(\IIO33.I2.net209 ), .d1(GND), .sl0(GND), .x(\IIO33.I2.net0153 ));
  invtd52_AVDD \IIO33.I2.I8  ( .a(\IIO33.I2.net0151 ), .en(VDD), .x(\LongBus_20<5> ));
  invtd52_AVDD \IIO33.I2.I26  ( .a(\IIO33.I2.net0153 ), .en(VDD), .x(\LongBus_21<13> ));
  buftd52C_UCCLAB \I1804.I38  ( .a(\LongBus_20<5> ), .en(VDD), .x(\net8311<10> ));
  buftd52C_UCCLAB \I1803.I30  ( .a(\LongBus_21<13> ), .en(VDD), .x(\net8320<2> ));
  buftd52C_UCCLAB \I3739.I38  ( .a(\net8311<10> ), .en(VDD), .x(\LongBus_79<5> ));
  buftd52C_UCCLAB \I3740.I30  ( .a(\net8320<2> ), .en(VDD), .x(\LongBus_78<13> ));
  buftd52_UCCLAB \ILAB0101.I4775.I38  ( .a(\LongBus_79<5> ), .en(VDD), .x(\LongBus_1<5> ));
  inv_4_UCCLAB \ILAB0102.ILE1605.I712  ( .a(\LongBus_1<5> ), .x(\ILAB0102.ILE1605.net0562 ));
  inv_4_UCCLAB \ILAB0101.ILE1613.I712  ( .a(\LongBus_1<5> ), .x(\ILAB0101.ILE1613.net0562 ));
  inv_4_UCCLAB \ILAB0101.ILE1516.I713  ( .a(\LongBus_78<13> ), .x(\ILAB0101.ILE1516.net01342 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1605.Iho3  ( .en(GND), .in(\ILAB0102.ILE1605.net0562 ), .out(\ILAB0102.net15864 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1303.Iho2  ( .en(GND), .in(\ILAB0101.ILE1516.net01342 ), .out(\ILAB0102.net16628 ));
  mux2i_P_UCCLAB \IIO33.I3.I25  ( .d0(\IIO33.I3.net209 ), .d1(GND), .sl0(GND), .x(\IIO33.I3.net0153 ));
  invtd52_AVDD \IIO33.I3.I26  ( .a(\IIO33.I3.net0153 ), .en(VDD), .x(\LongBus_21<12> ));
  buftd52C_UCCLAB \I1803.I33  ( .a(\LongBus_21<12> ), .en(VDD), .x(\net8320<3> ));
  inv_4_UCCLAB \ILAB0401.ILE0816.I715  ( .a(\net8320<3> ), .x(\ILAB0401.ILE0816.net01339 ));
  inv_8_UCCLAB \ILAB0401.ILE0816.I666  ( .a(\ILAB0401.ILE0816.net01339 ), .x(\net16243<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0812.Ihi7  ( .en(GND), .in(\ILAB0401.ILE0816.net01339 ), .out(\ILAB0401.net17977 ));
  buf4_12_UCCLAB \ILAB0401.I4373  ( .a(\net16243<1> ), .x(\ILAB0401.net27353 ));
  buftid52C_UCCLAB \ILAB0401.I4431  ( .a(\ILAB0401.net27353 ), .ne(GND), .x(\net8320<13> ));
  buftd52C_UCCLAB \I3740.I7  ( .a(\net8320<13> ), .en(VDD), .x(\LongBus_78<2> ));
  mux2i_P_UCCLAB \IIO10.I5.I16  ( .d0(\LongBus_78<2> ), .d1(GND), .sl0(GND), .x(\IIO10.I5.net197 ));
  mux2i_P_UCCLAB \IIO33.I4.I25  ( .d0(\IIO33.I4.net209 ), .d1(GND), .sl0(GND), .x(\IIO33.I4.net0153 ));
  invtd52_AVDD \IIO33.I4.I26  ( .a(\IIO33.I4.net0153 ), .en(VDD), .x(\LongBus_21<11> ));
  buftd52C_UCCLAB \I1803.I22  ( .a(\LongBus_21<11> ), .en(VDD), .x(\net8320<4> ));
  inv_4_UCCLAB \ILAB0401.ILE1016.I714  ( .a(\net8320<4> ), .x(\ILAB0401.ILE1016.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE1012.Ihi7  ( .en(GND), .in(\ILAB0401.ILE1016.net01345 ), .out(\ILAB0401.net24322 ));
  mux2i_P_UCCLAB \IIO33.I5.I25  ( .d0(\IIO33.I5.net209 ), .d1(GND), .sl0(GND), .x(\IIO33.I5.net0153 ));
  invtd52_AVDD \IIO33.I5.I26  ( .a(\IIO33.I5.net0153 ), .en(VDD), .x(\LongBus_21<10> ));
  buftd52_UCCLAB \ILAB1001.I4801.I25  ( .a(\LongBus_21<10> ), .en(VDD), .x(\LongBus_19<10> ));
  buftd52C_UCCLAB \I1803.I25  ( .a(\LongBus_21<10> ), .en(VDD), .x(\net8320<5> ));
  buftd52_UCCLAB \ILAB0401.I4773.I25  ( .a(\net8320<5> ), .en(VDD), .x(\LongBus_6<10> ));
  buftd52C_UCCLAB \I3740.I25  ( .a(\net8320<5> ), .en(VDD), .x(\LongBus_78<10> ));
  buftd52_UCCLAB \ILAB0402.I4772.I24  ( .a(\LongBus_6<10> ), .en(VDD), .x(\net8296<5> ));
  buftd52_UCCLAB \ILAB0402.I4773.I24  ( .a(\LongBus_6<10> ), .en(VDD), .x(\net8287<5> ));
  buftd52_UCCLAB \ILAB0201.I4773.I25  ( .a(\LongBus_78<10> ), .en(VDD), .x(\LongBus_2<10> ));
  buftd52_UCCLAB \ILAB0101.I4801.I25  ( .a(\LongBus_78<10> ), .en(VDD), .x(\LongBus_1<10> ));
  inv_4_UCCLAB \ILAB0401.ILE0716.I715  ( .a(\net8320<5> ), .x(\ILAB0401.ILE0716.net01339 ));
  buftd52C_UCCLAB \I3742.I25  ( .a(\net8287<5> ), .en(VDD), .x(\LongBus_72<10> ));
  buftd52C_UCCLAB \I3741.I25  ( .a(\net8296<5> ), .en(VDD), .x(\LongBus_73<10> ));
  inv_4_UCCLAB \ILAB0401.ILE0113.I715  ( .a(\LongBus_6<10> ), .x(\ILAB0401.ILE0113.net01339 ));
  inv_4_UCCLAB \ILAB0402.ILE0102.I715  ( .a(\LongBus_6<10> ), .x(\ILAB0402.ILE0102.net01339 ));
  inv_4_UCCLAB \ILAB1001.ILE1610.I712  ( .a(\LongBus_19<10> ), .x(\ILAB1001.ILE1610.net0562 ));
  inv_4_UCCLAB \ILAB0101.ILE0216.I715  ( .a(\LongBus_78<10> ), .x(\ILAB0101.ILE0216.net01339 ));
  inv_4_UCCLAB \ILAB0102.ILE1416.I715  ( .a(\LongBus_72<10> ), .x(\ILAB0102.ILE1416.net01339 ));
  inv_4_UCCLAB \ILAB0102.ILE0516.I715  ( .a(\LongBus_72<10> ), .x(\ILAB0102.ILE0516.net01339 ));
  inv_4_UCCLAB \ILAB0102.ILE0716.I715  ( .a(\LongBus_72<10> ), .x(\ILAB0102.ILE0716.net01339 ));
  inv_4_UCCLAB \ILAB0102.ILE0316.I715  ( .a(\LongBus_72<10> ), .x(\ILAB0102.ILE0316.net01339 ));
  inv_4_UCCLAB \ILAB0102.ILE1216.I715  ( .a(\LongBus_72<10> ), .x(\ILAB0102.ILE1216.net01339 ));
  inv_4_UCCLAB \ILAB0302.ILE1501.I715  ( .a(\LongBus_73<10> ), .x(\ILAB0302.ILE1501.net01339 ));
  inv_4_UCCLAB \ILAB0102.ILE0801.I715  ( .a(\LongBus_73<10> ), .x(\ILAB0102.ILE0801.net01339 ));
  inv_4_UCCLAB \ILAB0102.ILE0601.I715  ( .a(\LongBus_73<10> ), .x(\ILAB0102.ILE0601.net01339 ));
  inv_4_UCCLAB \ILAB0102.ILE0501.I715  ( .a(\LongBus_73<10> ), .x(\ILAB0102.ILE0501.net01339 ));
  inv_4_UCCLAB \ILAB0102.ILE0401.I715  ( .a(\LongBus_73<10> ), .x(\ILAB0102.ILE0401.net01339 ));
  inv_4_UCCLAB \ILAB0202.ILE0108.I715  ( .a(\LongBus_2<10> ), .x(\ILAB0202.ILE0108.net01339 ));
  inv_4_UCCLAB \ILAB0202.ILE0106.I715  ( .a(\LongBus_2<10> ), .x(\ILAB0202.ILE0106.net01339 ));
  inv_4_UCCLAB \ILAB0103.ILE1602.I711  ( .a(\LongBus_1<10> ), .x(\ILAB0103.ILE1602.net0560 ));
  inv_4_UCCLAB \ILAB0102.ILE1607.I712  ( .a(\LongBus_1<10> ), .x(\ILAB0102.ILE1607.net0562 ));
  inv_4_UCCLAB \ILAB0102.ILE1101.I715  ( .a(\LongBus_73<10> ), .x(\ILAB0102.ILE1101.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1201.Iho1  ( .en(GND), .in(\ILAB0102.ILE1216.net01339 ), .out(\ILAB0103.net15502 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0512.Ihi7  ( .en(GND), .in(\ILAB0102.ILE0516.net01339 ), .out(\ILAB0102.net19462 ));
  sw_b_v2_inv_UCCLAB \ILAB0101.ILE0216.Iho1  ( .en(GND), .in(\ILAB0101.ILE0216.net01339 ), .out(\net17230<6> ));
  mux2i_P_UCCLAB \IIO33.I5.I27  ( .d0(\IIO33.I5.net209 ), .d1(GND), .sl0(GND), .x(\IIO33.I5.net0151 ));
  invtd52_AVDD \IIO33.I5.I8  ( .a(\IIO33.I5.net0151 ), .en(VDD), .x(\LongBus_20<2> ));
  buftd52C_UCCLAB \I1804.I7  ( .a(\LongBus_20<2> ), .en(VDD), .x(\net8311<13> ));
  buftd52_UCCLAB \ILAB0401.I4772.I7  ( .a(\net8311<13> ), .en(VDD), .x(\LongBus_6<2> ));
  buftd52_UCCLAB \ILAB0403.I4772.I6  ( .a(\LongBus_6<2> ), .en(VDD), .x(\net8299<13> ));
  buftd52C_UCCLAB \I3743.I7  ( .a(\net8299<13> ), .en(VDD), .x(\LongBus_71<2> ));
  inv_4_UCCLAB \ILAB0401.ILE0816.I713  ( .a(\net8320<5> ), .x(\ILAB0401.ILE0816.net01342 ));
  inv_4_UCCLAB \ILAB0201.ILE0316.I714  ( .a(\LongBus_78<10> ), .x(\ILAB0201.ILE0316.net01345 ));
  inv_4_UCCLAB \ILAB0102.ILE1608.I712  ( .a(\LongBus_1<10> ), .x(\ILAB0102.ILE1608.net0562 ));
  inv_4_UCCLAB \ILAB0103.ILE0401.I715  ( .a(\LongBus_71<2> ), .x(\ILAB0103.ILE0401.net01339 ));
  inv_4_UCCLAB \ILAB0103.ILE0701.I715  ( .a(\LongBus_71<2> ), .x(\ILAB0103.ILE0701.net01339 ));
  inv_4_UCCLAB \ILAB0103.ILE0201.I715  ( .a(\LongBus_71<2> ), .x(\ILAB0103.ILE0201.net01339 ));
  inv_4_UCCLAB \ILAB0102.ILE1301.I713  ( .a(\LongBus_73<10> ), .x(\ILAB0102.ILE1301.net01342 ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0102.Ivo3  ( .en(GND), .in(\ILAB0402.ILE0102.net01339 ), .out(\ILAB0402.net26775 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0712.Ihi7  ( .en(GND), .in(\ILAB0401.ILE0716.net01339 ), .out(\ILAB0401.net21037 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1213.Ihi7  ( .en(GND), .in(\ILAB0102.ILE1216.net01339 ), .out(\ILAB0102.net16267 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0516.Iho1  ( .en(GND), .in(\ILAB0102.ILE0516.net01339 ), .out(\net10423<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0214.Ihi7  ( .en(GND), .in(\ILAB0103.ILE0201.net01339 ), .out(\ILAB0102.net25537 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0202.Iho1  ( .en(GND), .in(\ILAB0103.ILE0201.net01339 ), .out(\ILAB0103.net26752 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0401.Ivo3  ( .en(GND), .in(\ILAB0103.ILE0401.net01339 ), .out(\ILAB0103.net20655 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0504.Iho1  ( .en(GND), .in(\net10423<6> ), .out(\ILAB0103.net24997 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0416.Iho2  ( .en(GND), .in(\ILAB0103.ILE0401.net01339 ), .out(\net10427<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1208.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1608.net0562 ), .out(\ILAB0102.net22639 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0602.Iho1  ( .en(GND), .in(\ILAB0102.ILE0601.net01339 ), .out(\ILAB0102.net26392 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0402.Iho3  ( .en(GND), .in(\net10427<5> ), .out(\ILAB0103.net26214 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1407.Ivi6  ( .en(GND), .in(\ILAB0102.ILE1607.net0562 ), .out(\ILAB0102.net25744 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0808.Ivi7  ( .en(GND), .in(\ILAB0102.net22639 ), .out(\ILAB0102.net18004 ));
  inv_4_UCCLAB \ILAB0401.ILE0316.I713  ( .a(\net8320<5> ), .x(\ILAB0401.ILE0316.net01342 ));
  inv_4_UCCLAB \ILAB0101.ILE0416.I713  ( .a(\LongBus_78<10> ), .x(\ILAB0101.ILE0416.net01342 ));
  inv_4_UCCLAB \ILAB0102.ILE1001.I714  ( .a(\LongBus_73<10> ), .x(\ILAB0102.ILE1001.net01345 ));
  inv_4_UCCLAB \ILAB0102.ILE1501.I715  ( .a(\LongBus_73<10> ), .x(\ILAB0102.ILE1501.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0301.ILE1513.Ivi6  ( .en(GND), .in(\ILAB0401.ILE0113.net01339 ), .out(\net16377<4> ));
  sw_b_v2_inv_UCCLAB \ILAB0301.ILE1613.Ivo1  ( .en(GND), .in(\net16377<4> ), .out(\net16279<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0101.ILE0816.Iho2  ( .en(GND), .in(\ILAB0102.ILE0801.net01339 ), .out(\net17206<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0401.Iho1  ( .en(GND), .in(\ILAB0101.ILE0416.net01342 ), .out(\ILAB0102.net20722 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0802.Iho3  ( .en(GND), .in(\net17206<5> ), .out(\ILAB0102.net26124 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0314.Ihi6  ( .en(GND), .in(\ILAB0401.ILE0316.net01342 ), .out(\ILAB0401.net23377 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0404.Iho2  ( .en(GND), .in(\ILAB0102.net20722 ), .out(\ILAB0102.net15548 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0305.Iho1  ( .en(GND), .in(\ILAB0102.ILE0601.net01339 ), .out(\ILAB0102.net23332 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1213.Ivi5  ( .en(GND), .in(\ILAB0102.ILE1216.net01339 ), .out(\ILAB0102.net21107 ));
  inv_8_UCCLAB \ILAB0103.ILE1602.I666  ( .a(\ILAB0103.ILE1602.net0560 ), .x(\ILAB0103.net20561 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0606.Iho1  ( .en(GND), .in(\ILAB0102.net26392 ), .out(\ILAB0102.net18562 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1107.Ivi7  ( .en(GND), .in(\ILAB0102.net25744 ), .out(\ILAB0102.net17194 ));
  buftd4_UCCLAB \ILAB0103.I231  ( .a(\ILAB0103.net20561 ), .en(VDD), .x(\ILAB0103.net027166 ));
  mux2p_2_UCCLAB \ILAB0103.I5605.I4  ( .d0(\ILAB0103.net027166 ), .d1(GND), .s0(GND), .x(\ILAB0103.I5605.net25 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1013.Ivi6  ( .en(GND), .in(\ILAB0102.net21107 ), .out(\ILAB0102.net21559 ));
  invd16_seth_UCCLAB \ILAB0103.I5605.I5  ( .a(\ILAB0103.I5605.net25 ), .c(VDD), .x(\ILAB0103.Clk_int<1> ));
  mux2d1i_1_P_UCCLAB \ILAB0103.I5366.I79  ( .d0(\ILAB0103.Clk_int<1> ), .d1i(GND), .sl0(GND), .x(\ILAB0103.I5366.net0110 ));
  invd52_UCCLAB \ILAB0103.I5366.I75  ( .a(\ILAB0103.I5366.net0110 ), .x(\ILAB0103.net15299<2> ));
  invd32_UCCLAB \ILAB0103.I5591.I2  ( .a(\ILAB0103.net15299<2> ), .x(\ILAB0103.Clk_LAB<1> ));
  inv_4_UCCLAB \ILAB0401.ILE0916.I715  ( .a(\net8320<5> ), .x(\ILAB0401.ILE0916.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0702.Iho1  ( .en(GND), .in(\ILAB0103.ILE0701.net01339 ), .out(\ILAB0103.net26437 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0604.Iho2  ( .en(GND), .in(\ILAB0102.ILE0801.net01339 ), .out(\ILAB0102.net25988 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0912.Ivo3  ( .en(GND), .in(\ILAB0102.ILE0716.net01339 ), .out(\ILAB0102.net21690 ));
  mux2i_P_UCCLAB \IIO33.I6.I25  ( .d0(\IIO33.I6.net209 ), .d1(GND), .sl0(GND), .x(\IIO33.I6.net0153 ));
  invtd52_AVDD \IIO33.I6.I26  ( .a(\IIO33.I6.net0153 ), .en(VDD), .x(\LongBus_21<9> ));
  buftd52C_UCCLAB \I1803.I21  ( .a(\LongBus_21<9> ), .en(VDD), .x(\net8320<6> ));
  buftd52C_UCCLAB \I3740.I21  ( .a(\net8320<6> ), .en(VDD), .x(\LongBus_78<9> ));
  inv_4_UCCLAB \ILAB0401.ILE1616.I714  ( .a(\net8320<6> ), .x(\ILAB0401.ILE1616.net01345 ));
  inv_4_UCCLAB \ILAB0201.ILE0316.I715  ( .a(\LongBus_78<9> ), .x(\ILAB0201.ILE0316.net01339 ));
  inv_8_UCCLAB \ILAB0201.ILE0316.I666  ( .a(\ILAB0201.ILE0316.net01339 ), .x(\net18362<1> ));
  buf4_12_UCCLAB \ILAB0201.I4398  ( .a(\net18362<1> ), .x(\ILAB0201.net27303 ));
  inv_8_UCCLAB \ILAB0401.ILE1616.I666  ( .a(\ILAB0401.ILE1616.net01345 ), .x(\net16235<1> ));
  buftid52C_UCCLAB \ILAB0201.I4420  ( .a(\ILAB0201.net27303 ), .ne(GND), .x(\LongBus_78<5> ));
  mux2i_P_UCCLAB \IIO10.I2.I16  ( .d0(\LongBus_78<5> ), .d1(GND), .sl0(GND), .x(\IIO10.I2.net197 ));
  buftd4_UCCLAB \ILAB0401.I178  ( .a(\net16235<1> ), .en(VDD), .x(\ILAB0401.net015238 ));
  mux2p_2_UCCLAB \ILAB0401.I5605.I2  ( .d0(GND), .d1(\ILAB0401.net015238 ), .s0(VDD), .x(\ILAB0401.I5605.net33 ));
  invd16_seth_UCCLAB \ILAB0401.I5605.I3  ( .a(\ILAB0401.I5605.net33 ), .c(VDD), .x(\ILAB0401.Clk_int<2> ));
  mux2d1i_1_P_UCCLAB \ILAB0401.I5366.I80  ( .d0(\ILAB0401.Clk_int<2> ), .d1i(GND), .sl0(GND), .x(\ILAB0401.I5366.net0106 ));
  invd52_UCCLAB \ILAB0401.I5366.I76  ( .a(\ILAB0401.I5366.net0106 ), .x(\ILAB0401.net15299<1> ));
  invd32_UCCLAB \ILAB0401.I5591.I1  ( .a(\ILAB0401.net15299<1> ), .x(\ILAB0401.Clk_LAB<2> ));
  sw_b_v2_inv_UCCLAB \ILAB0101.ILE0916.Iho3  ( .en(GND), .in(\ILAB0101.ILE0916.net2656 ), .out(\net17202<4> ));
  inv_8_UCCLAB \ILAB0101.ILE0916.I666  ( .a(\ILAB0101.ILE0916.net0541 ), .x(\net17148<1> ));
  buf4_12_UCCLAB \ILAB0101.I4401  ( .a(\net17148<1> ), .x(\ILAB0101.net27297 ));
  buftid52C_UCCLAB \ILAB0101.I4464  ( .a(\ILAB0101.net27297 ), .ne(GND), .x(\LongBus_78<6> ));
  mux2i_P_UCCLAB \IIO10.I1.I16  ( .d0(\LongBus_78<6> ), .d1(GND), .sl0(GND), .x(\IIO10.I1.net197 ));
  inv_8_UCCLAB \ILAB0101.ILE0215.I666  ( .a(\ILAB0101.ILE0215.net0541 ), .x(\ILAB0101.net23756 ));
  inv_8_UCCLAB \ILAB0101.ILE0216.I666  ( .a(\ILAB0101.net23756 ), .x(\net17155<1> ));
  buf4_12_UCCLAB \ILAB0101.I4402  ( .a(\net17155<1> ), .x(\ILAB0101.net27295 ));
  buftid52C_UCCLAB \ILAB0101.I4432  ( .a(\ILAB0101.net27295 ), .ne(GND), .x(\LongBus_78<4> ));
  mux2i_P_UCCLAB \IIO10.I3.I16  ( .d0(\LongBus_78<4> ), .d1(GND), .sl0(GND), .x(\IIO10.I3.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB1001.ILE1410.Ihi7  ( .en(GND), .in(\ILAB1001.ILE1410.net2656 ), .out(\ILAB1001.net21127 ));
  sw_b_v2_inv_UCCLAB \ILAB1001.ILE1410.Iho1  ( .en(GND), .in(\ILAB1001.ILE1410.net2656 ), .out(\ILAB1001.net24007 ));
  sw_b_v2_inv_UCCLAB \ILAB1001.ILE1406.Ihi7  ( .en(GND), .in(\ILAB1001.net21127 ), .out(\ILAB1001.net26302 ));
  sw_b_v2_inv_UCCLAB \ILAB1001.ILE1414.Iho1  ( .en(GND), .in(\ILAB1001.net24007 ), .out(\net16578<1> ));
  inv_8_UCCLAB \ILAB1001.ILE1416.I666  ( .a(\net16578<1> ), .x(\net16539<1> ));
  buf4_12_UCCLAB \ILAB1001.I4369  ( .a(\net16539<1> ), .x(\ILAB1001.net27361 ));
  inv_8_UCCLAB \ILAB1001.ILE1602.I666  ( .a(\ILAB1001.net26302 ), .x(\ILAB1001.net20561 ));
  buftd4_UCCLAB \ILAB1001.I231  ( .a(\ILAB1001.net20561 ), .en(VDD), .x(\ILAB1001.net027166 ));
  buftd4_UCCLAB \ILAB1001.I233  ( .a(\ILAB1001.net20561 ), .en(VDD), .x(\ILAB1001.net027160 ));
  mux2p_2_UCCLAB \ILAB1001.I5605.I4  ( .d0(\ILAB1001.net027166 ), .d1(GND), .s0(GND), .x(\ILAB1001.I5605.net25 ));
  mux2p_2_UCCLAB \ILAB1001.I5605.I7  ( .d0(\ILAB1001.net027160 ), .d1(GND), .s0(GND), .x(\ILAB1001.I5605.net21 ));
  invd16_seth_UCCLAB \ILAB1001.I5605.I6  ( .a(\ILAB1001.I5605.net21 ), .c(VDD), .x(\ILAB1001.Clk_int<0> ));
  invd16_seth_UCCLAB \ILAB1001.I5605.I5  ( .a(\ILAB1001.I5605.net25 ), .c(VDD), .x(\ILAB1001.Clk_int<1> ));
  mux2p_2_UCCLAB \ILAB1001.I5366.I82  ( .d0(\ILAB1001.Clk_int<0> ), .d1(GND), .s0(GND), .x(\ILAB1001.I5366.net0119 ));
  mux2p_2_UCCLAB \ILAB1001.I5366.I83  ( .d0(\ILAB1001.Clk_int<1> ), .d1(GND), .s0(GND), .x(\ILAB1001.I5366.net0122 ));
  invtd56_clk_UCCLAB \ILAB1001.I5366.I6  ( .a(\ILAB1001.I5366.net0119 ), .en(VDD), .x(\net16523<1> ));
  invtd56_clk_UCCLAB \ILAB1001.I5366.I8  ( .a(\ILAB1001.I5366.net0122 ), .en(VDD), .x(\net16523<0> ));
  invtd56_UCCLAB \I3706.I4  ( .a(\net16523<1> ), .en(VDD), .x(\net10305<1> ));
  invtd56_UCCLAB \I3706.I3  ( .a(\net16523<0> ), .en(VDD), .x(\net10305<0> ));
  mux2_1_clk_P_UCCLAB \I3590.I21  ( .d0(\net10305<1> ), .d1(GND), .sl0(GND), .x(\I3590.net052 ));
  mux2_1_clk_P_UCCLAB \I3590.I16  ( .d0(\net10305<0> ), .d1(GND), .sl0(GND), .x(\I3590.net073 ));
  mux2_1_clk_P_UCCLAB \I3590.I20  ( .d0(\net10305<0> ), .d1(GND), .sl0(GND), .x(\I3590.net059 ));
  mux4p_0_UCCLAB \I3590.I12  ( .d0(GND), .d1(GND), .d2(GND), .d3(\I3590.net073 ), .sl0(VDD), .sl1(VDD), .x(\I3590.net84 ));
  mux4p_0_UCCLAB \I3590.I14  ( .d0(GND), .d1(GND), .d2(GND), .d3(\I3590.net059 ), .sl0(VDD), .sl1(VDD), .x(\I3590.net72 ));
  mux4p_0_UCCLAB \I3590.I15  ( .d0(GND), .d1(GND), .d2(GND), .d3(\I3590.net052 ), .sl0(VDD), .sl1(VDD), .x(\I3590.net66 ));
  invtd56_pd_clk_UCCLAB \I3590.I0  ( .a(\I3590.net84 ), .en(VDD), .x(\net10262<0> ));
  invtd56_pd_clk_UCCLAB \I3590.I7  ( .a(\I3590.net72 ), .en(VDD), .x(\net10262<2> ));
  invtd56_pd_clk_UCCLAB \I3590.I9  ( .a(\I3590.net66 ), .en(VDD), .x(\net10262<3> ));
  mux2p_2_UCCLAB \I3689.I3  ( .d0(\net10262<2> ), .d1(GND), .s0(GND), .x(\I3689.net39 ));
  mux2p_2_UCCLAB \I3690.I6  ( .d0(\net10262<0> ), .d1(GND), .s0(GND), .x(\I3690.net47 ));
  mux2p_2_UCCLAB \I3689.I2  ( .d0(\net10262<3> ), .d1(GND), .s0(GND), .x(\I3689.net35 ));
  invtd56_pd_clk_UCCLAB \I3689.I7  ( .a(\I3689.net39 ), .en(VDD), .x(\net20977<2> ));
  invtd56_pd_clk_UCCLAB \I3690.I0  ( .a(\I3690.net47 ), .en(VDD), .x(\net20974<0> ));
  invtd56_pd_clk_UCCLAB \I3689.I9  ( .a(\I3689.net35 ), .en(VDD), .x(\net20977<3> ));
  buftid52C_UCCLAB \ILAB1001.I4419  ( .a(\ILAB1001.net27361 ), .ne(GND), .x(\LongBus_21<3> ));
  invtd56_pd_clk_UCCLAB \I3648.I3  ( .a(\net20977<2> ), .en(VDD), .x(\net16222<2> ));
  invtd56_pd_clk_UCCLAB \I3648.I4  ( .a(\net20977<3> ), .en(VDD), .x(\net16222<3> ));
  buftd52C_UCCLAB \I1803.I9  ( .a(\LongBus_21<3> ), .en(VDD), .x(\net8320<12> ));
  nand2_1_UCCLAB \ILAB0402.I5366.I71  ( .a(VDD), .b(\net16222<2> ), .x(\ILAB0402.I5366.net70 ));
  nand2_1_UCCLAB \ILAB0302.I5366.I71  ( .a(VDD), .b(\net16222<2> ), .x(\ILAB0302.I5366.net70 ));
  nand2_1_UCCLAB \ILAB0401.I5366.I0  ( .a(VDD), .b(\net16222<3> ), .x(\ILAB0401.I5366.net64 ));
  buftd52C_UCCLAB \I3740.I9  ( .a(\net8320<12> ), .en(VDD), .x(\LongBus_78<3> ));
  mux2d1i_1_P_UCCLAB \ILAB0302.I5366.I79  ( .d0(GND), .d1i(\ILAB0302.I5366.net70 ), .sl0(VDD), .x(\ILAB0302.I5366.net0110 ));
  mux2d1i_1_P_UCCLAB \ILAB0401.I5366.I78  ( .d0(GND), .d1i(\ILAB0401.I5366.net64 ), .sl0(VDD), .x(\ILAB0401.I5366.net0114 ));
  mux2d1i_1_P_UCCLAB \ILAB0402.I5366.I79  ( .d0(GND), .d1i(\ILAB0402.I5366.net70 ), .sl0(VDD), .x(\ILAB0402.I5366.net0110 ));
  mux2i_P_UCCLAB \IIO10.I4.I16  ( .d0(\LongBus_78<3> ), .d1(GND), .sl0(GND), .x(\IIO10.I4.net197 ));
  invd52_UCCLAB \ILAB0402.I5366.I75  ( .a(\ILAB0402.I5366.net0110 ), .x(\ILAB0402.net15299<2> ));
  invd52_UCCLAB \ILAB0302.I5366.I75  ( .a(\ILAB0302.I5366.net0110 ), .x(\ILAB0302.net15299<2> ));
  invd52_UCCLAB \ILAB0401.I5366.I74  ( .a(\ILAB0401.I5366.net0114 ), .x(\ILAB0401.net15299<3> ));
  invd32_UCCLAB \ILAB0402.I5591.I2  ( .a(\ILAB0402.net15299<2> ), .x(\ILAB0402.Clk_LAB<1> ));
  invd32_UCCLAB \ILAB0302.I5591.I2  ( .a(\ILAB0302.net15299<2> ), .x(\ILAB0302.Clk_LAB<1> ));
  invd32_UCCLAB \ILAB0401.I5591.I3  ( .a(\ILAB0401.net15299<3> ), .x(\ILAB0401.Clk_LAB<0> ));
  mux2p_2_UCCLAB \I3690.I2  ( .d0(\net10262<3> ), .d1(GND), .s0(GND), .x(\I3690.net35 ));
  invtd56_pd_clk_UCCLAB \I3690.I9  ( .a(\I3690.net35 ), .en(VDD), .x(\net20974<3> ));
  invtd56_pd_clk_UCCLAB \I3651.I4  ( .a(\net20974<3> ), .en(VDD), .x(\GCLK_s1<0> ));
  invtd56_pd_clk_UCCLAB \I3652.I1  ( .a(\net20974<0> ), .en(VDD), .x(\net20955<0> ));
  nand2_1_UCCLAB \ILAB0103.I5366.I73  ( .a(VDD), .b(\net20955<0> ), .x(\ILAB0103.I5366.net66 ));
  nand2_1_UCCLAB \ILAB0201.I5366.I0  ( .a(VDD), .b(\GCLK_s1<0> ), .x(\ILAB0201.I5366.net64 ));
  nand2_1_UCCLAB \ILAB0101.I5366.I0  ( .a(VDD), .b(\GCLK_s1<0> ), .x(\ILAB0101.I5366.net64 ));
  nand2_1_UCCLAB \ILAB0102.I5366.I0  ( .a(VDD), .b(\GCLK_s1<0> ), .x(\ILAB0102.I5366.net64 ));
  mux2d1i_1_P_UCCLAB \ILAB0103.I5366.I81  ( .d0(GND), .d1i(\ILAB0103.I5366.net66 ), .sl0(VDD), .x(\ILAB0103.I5366.net0102 ));
  mux2d1i_1_P_UCCLAB \ILAB0201.I5366.I78  ( .d0(GND), .d1i(\ILAB0201.I5366.net64 ), .sl0(VDD), .x(\ILAB0201.I5366.net0114 ));
  mux2d1i_1_P_UCCLAB \ILAB0101.I5366.I78  ( .d0(GND), .d1i(\ILAB0101.I5366.net64 ), .sl0(VDD), .x(\ILAB0101.I5366.net0114 ));
  mux2d1i_1_P_UCCLAB \ILAB0102.I5366.I78  ( .d0(GND), .d1i(\ILAB0102.I5366.net64 ), .sl0(VDD), .x(\ILAB0102.I5366.net0114 ));
  invd52_UCCLAB \ILAB0101.I5366.I74  ( .a(\ILAB0101.I5366.net0114 ), .x(\ILAB0101.net15299<3> ));
  invd52_UCCLAB \ILAB0201.I5366.I74  ( .a(\ILAB0201.I5366.net0114 ), .x(\ILAB0201.net15299<3> ));
  invd52_UCCLAB \ILAB0103.I5366.I77  ( .a(\ILAB0103.I5366.net0102 ), .x(\ILAB0103.net15299<0> ));
  invd52_UCCLAB \ILAB0102.I5366.I74  ( .a(\ILAB0102.I5366.net0114 ), .x(\ILAB0102.net15299<3> ));
  invd32_UCCLAB \ILAB0101.I5591.I3  ( .a(\ILAB0101.net15299<3> ), .x(\ILAB0101.Clk_LAB<0> ));
  invd32_UCCLAB \ILAB0201.I5591.I3  ( .a(\ILAB0201.net15299<3> ), .x(\ILAB0201.Clk_LAB<0> ));
  invd32_UCCLAB \ILAB0102.I5591.I3  ( .a(\ILAB0102.net15299<3> ), .x(\ILAB0102.Clk_LAB<0> ));
  invd32_UCCLAB \ILAB0103.I5591.I0  ( .a(\ILAB0103.net15299<0> ), .x(\ILAB0103.Clk_LAB<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0403.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0403.net2656 ), .out(\net10430<6> ));
  inv_8_UCCLAB \ILAB0102.ILE0103.I666  ( .a(\net10430<6> ), .x(\ILAB0102.net26726 ));
  buf4_12_UCCLAB \ILAB0102.I4362  ( .a(\ILAB0102.net26726 ), .x(\ILAB0102.net40017 ));
  buftd52C_UCCLAB \ILAB0102.I4442  ( .a(\ILAB0102.net40017 ), .en(VDD), .x(\LongBus_0<1> ));
  buftd52_UCCLAB \ILAB0101.I4773.I4  ( .a(\LongBus_0<1> ), .en(VDD), .x(\LongBus_78<1> ));
  mux2i_P_UCCLAB \IIO10.I6.I16  ( .d0(\LongBus_78<1> ), .d1(GND), .sl0(GND), .x(\IIO10.I6.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0403.Ivo2  ( .en(GND), .in(\ILAB0102.ILE0403.net2656 ), .out(\ILAB0102.net17687 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0404.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0404.net2656 ), .out(\net10426<6> ));
  inv_8_UCCLAB \ILAB0102.ILE0104.I666  ( .a(\net10426<6> ), .x(\ILAB0102.net22856 ));
  buf4_12_UCCLAB \ILAB0102.I4378  ( .a(\ILAB0102.net22856 ), .x(\ILAB0102.net37425 ));
  buftd52C_UCCLAB \ILAB0102.I4435  ( .a(\ILAB0102.net37425 ), .en(VDD), .x(\LongBus_0<0> ));
  buftd52_UCCLAB \ILAB0101.I4773.I1  ( .a(\LongBus_0<0> ), .en(VDD), .x(\LongBus_78<0> ));
  mux2i_P_UCCLAB \IIO10.I7.I16  ( .d0(\LongBus_78<0> ), .d1(GND), .sl0(GND), .x(\IIO10.I7.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0404.Ivo3  ( .en(GND), .in(\ILAB0102.ILE0404.net2656 ), .out(\ILAB0102.net25020 ));
  inv_8_UCCLAB \ILAB0102.ILE0801.I666  ( .a(\ILAB0102.ILE0801.net0541 ), .x(\net17149<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0801.Ivi6  ( .en(GND), .in(\ILAB0102.ILE0801.net2656 ), .out(\ILAB0102.net20929 ));
  buf4_12_UCCLAB \ILAB0102.I4374  ( .a(\net17149<0> ), .x(\ILAB0102.net39222 ));
  buftid52C_UCCLAB \ILAB0102.I4476  ( .a(\ILAB0102.net39222 ), .ne(GND), .x(\LongBus_73<15> ));
  mux2i_P_UCCLAB \IIO11.I0.I16  ( .d0(GND), .d1(\LongBus_73<15> ), .sl0(VDD), .x(\IIO11.I0.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0801.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0801.net2656 ), .out(\ILAB0102.net20704 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0801.Iho2  ( .en(GND), .in(\ILAB0102.ILE0801.net2656 ), .out(\ILAB0102.net20678 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0601.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0601.net2656 ), .out(\ILAB0102.net20614 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0601.Iho2  ( .en(GND), .in(\ILAB0102.ILE0601.net2656 ), .out(\ILAB0102.net20588 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0601.Ivi5  ( .en(GND), .in(\ILAB0102.ILE0601.net2656 ), .out(\ILAB0102.net20612 ));
  inv_8_UCCLAB \ILAB0102.ILE0601.I666  ( .a(\ILAB0102.ILE0601.net0541 ), .x(\net17151<0> ));
  buf4_12_UCCLAB \ILAB0102.I4412  ( .a(\net17151<0> ), .x(\ILAB0102.net38382 ));
  buftid52C_UCCLAB \ILAB0102.I4456  ( .a(\ILAB0102.net38382 ), .ne(GND), .x(\LongBus_73<14> ));
  mux2i_P_UCCLAB \IIO11.I1.I16  ( .d0(GND), .d1(\LongBus_73<14> ), .sl0(VDD), .x(\IIO11.I1.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0605.Ihi5  ( .en(GND), .in(\ILAB0102.ILE0605.net2656 ), .out(\ILAB0102.net17663 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0605.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0605.net2656 ), .out(\ILAB0102.net15799 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0303.Ihi6  ( .en(GND), .in(\ILAB0102.net15799 ), .out(\net17226<6> ));
  inv_8_UCCLAB \ILAB0102.ILE0301.I666  ( .a(\net17226<6> ), .x(\net17154<0> ));
  buf4_12_UCCLAB \ILAB0102.I4394  ( .a(\net17154<0> ), .x(\ILAB0102.net38964 ));
  buftid52C_UCCLAB \ILAB0102.I4454  ( .a(\ILAB0102.net38964 ), .ne(GND), .x(\LongBus_73<13> ));
  mux2i_P_UCCLAB \IIO11.I2.I16  ( .d0(GND), .d1(\LongBus_73<13> ), .sl0(VDD), .x(\IIO11.I2.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0606.Ivo1  ( .en(GND), .in(\ILAB0102.ILE0606.net2656 ), .out(\ILAB0102.net18229 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0606.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0606.net2656 ), .out(\ILAB0102.net18589 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0703.Ihi7  ( .en(GND), .in(\ILAB0102.net18229 ), .out(\net17210<3> ));
  inv_8_UCCLAB \ILAB0102.ILE0701.I666  ( .a(\net17210<3> ), .x(\net17150<0> ));
  buf4_12_UCCLAB \ILAB0102.I4395  ( .a(\net17150<0> ), .x(\ILAB0102.net39618 ));
  buftid52C_UCCLAB \ILAB0102.I4455  ( .a(\ILAB0102.net39618 ), .ne(GND), .x(\LongBus_73<12> ));
  mux2i_P_UCCLAB \IIO11.I3.I16  ( .d0(GND), .d1(\LongBus_73<12> ), .sl0(VDD), .x(\IIO11.I3.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0508.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0508.net2656 ), .out(\Fast_out_28<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0508.Ihi7  ( .en(GND), .in(\ILAB0102.ILE0508.net2656 ), .out(\ILAB0102.net24997 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0504.Ihi7  ( .en(GND), .in(\ILAB0102.net24997 ), .out(\net17218<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0508.Ivo3  ( .en(GND), .in(\ILAB0102.ILE0508.net2656 ), .out(\ILAB0102.net19620 ));
  inv_8_UCCLAB \ILAB0102.ILE0501.I666  ( .a(\net17218<6> ), .x(\net17152<0> ));
  buf4_12_UCCLAB \ILAB0102.I4367  ( .a(\net17152<0> ), .x(\ILAB0102.net39858 ));
  buftid52C_UCCLAB \ILAB0102.I4470  ( .a(\ILAB0102.net39858 ), .ne(GND), .x(\LongBus_73<11> ));
  mux2i_P_UCCLAB \IIO11.I4.I16  ( .d0(GND), .d1(\LongBus_73<11> ), .sl0(VDD), .x(\IIO11.I4.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0610.Ivo3  ( .en(GND), .in(\ILAB0102.ILE0610.net2656 ), .out(\ILAB0102.net24165 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0610.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0610.net2656 ), .out(\ILAB0102.net24124 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0210.Ivi7  ( .en(GND), .in(\ILAB0102.net24124 ), .out(\ELLR9_28<5> ));
  inv_8_UCCLAB \ILAB0102.ILE0110.I666  ( .a(\ELLR9_28<5> ), .x(\ILAB0102.net16421 ));
  buf4_12_UCCLAB \ILAB0102.I4363  ( .a(\ILAB0102.net16421 ), .x(\ILAB0102.net40197 ));
  buftd52C_UCCLAB \ILAB0102.I4437  ( .a(\ILAB0102.net40197 ), .en(VDD), .x(\LongBus_0<2> ));
  buftd52_UCCLAB \ILAB0102.I4773.I6  ( .a(\LongBus_0<2> ), .en(VDD), .x(\LongBus_72<2> ));
  mux2i_P_UCCLAB \IIO11.I5.I16  ( .d0(\LongBus_72<2> ), .d1(GND), .sl0(GND), .x(\IIO11.I5.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1012.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1012.net2656 ), .out(\ILAB0102.net21694 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1012.Ivi5  ( .en(GND), .in(\ILAB0102.ILE1012.net2656 ), .out(\ILAB0102.net21692 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1012.Ivo1  ( .en(GND), .in(\ILAB0102.ILE1012.net2656 ), .out(\ILAB0102.net19399 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0812.Ivi6  ( .en(GND), .in(\ILAB0102.net21692 ), .out(\ILAB0102.net18949 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1412.Ivo1  ( .en(GND), .in(\ILAB0102.net19399 ), .out(\net18548<1> ));
  inv_8_UCCLAB \ILAB0202.ILE0112.I666  ( .a(\net18548<1> ), .x(\ILAB0202.net23216 ));
  buf4_12_UCCLAB \ILAB0202.I4371  ( .a(\ILAB0202.net23216 ), .x(\ILAB0202.net40041 ));
  buftd52C_UCCLAB \ILAB0202.I4436  ( .a(\ILAB0202.net40041 ), .en(VDD), .x(\LongBus_2<9> ));
  buftd52_UCCLAB \ILAB0202.I4772.I20  ( .a(\LongBus_2<9> ), .en(VDD), .x(\LongBus_73<9> ));
  mux2i_P_UCCLAB \IIO11.I6.I16  ( .d0(GND), .d1(\LongBus_73<9> ), .sl0(VDD), .x(\IIO11.I6.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1012.Ihi5  ( .en(GND), .in(\ILAB0102.ILE1012.net2656 ), .out(\ILAB0102.net24863 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1307.Ihi5  ( .en(GND), .in(\ILAB0102.ILE1307.net2656 ), .out(\ILAB0102.net15908 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1307.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1307.net2656 ), .out(\ILAB0102.net17149 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0907.Ivi7  ( .en(GND), .in(\ILAB0102.net17149 ), .out(\ILAB0102.net25969 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1307.Ivo1  ( .en(GND), .in(\ILAB0102.ILE1307.net2656 ), .out(\net18568<0> ));
  inv_8_UCCLAB \ILAB0102.ILE1607.I666  ( .a(\net18568<0> ), .x(\ILAB0102.net18266 ));
  buf4_12_UCCLAB \ILAB0102.I4357  ( .a(\ILAB0102.net18266 ), .x(\ILAB0102.net38148 ));
  buftd52C_UCCLAB \ILAB0102.I4425  ( .a(\ILAB0102.net38148 ), .en(VDD), .x(\LongBus_1<8> ));
  buftd52_UCCLAB \ILAB0102.I4775.I19  ( .a(\LongBus_1<8> ), .en(VDD), .x(\LongBus_73<8> ));
  mux2i_P_UCCLAB \IIO11.I7.I16  ( .d0(GND), .d1(\LongBus_73<8> ), .sl0(VDD), .x(\IIO11.I7.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1212.Ivo1  ( .en(GND), .in(\ILAB0102.ILE1212.net2656 ), .out(\net10337<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1212.Ivi5  ( .en(GND), .in(\ILAB0102.ILE1212.net2656 ), .out(\ILAB0102.net21377 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1012.Ivi6  ( .en(GND), .in(\ILAB0102.net21377 ), .out(\ILAB0102.net21784 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0712.Ivi7  ( .en(GND), .in(\ILAB0102.net21784 ), .out(\ILAB0102.net19939 ));
  inv_8_UCCLAB \ILAB0102.ILE1612.I666  ( .a(\net10337<3> ), .x(\ILAB0102.net22001 ));
  buf4_12_UCCLAB \ILAB0102.I4365  ( .a(\ILAB0102.net22001 ), .x(\ILAB0102.net39579 ));
  buftd52C_UCCLAB \ILAB0102.I4424  ( .a(\ILAB0102.net39579 ), .en(VDD), .x(\LongBus_1<7> ));
  buftd52_UCCLAB \ILAB0103.I4801.I36  ( .a(\LongBus_1<7> ), .en(VDD), .x(\LongBus_70<7> ));
  mux2i_P_UCCLAB \IIO12.I0.I16  ( .d0(\LongBus_70<7> ), .d1(GND), .sl0(GND), .x(\IIO12.I0.net197 ));
  inv_8_UCCLAB \ILAB0102.ILE0714.I666  ( .a(\ILAB0102.ILE0714.net0541 ), .x(\ILAB0102.net19976 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0714.Iho2  ( .en(GND), .in(\ILAB0102.ILE0714.net2656 ), .out(\ILAB0102.net22388 ));
  inv_4_UCCLAB \ILAB0102.ILE0613.I710  ( .a(\ILAB0102.net19976 ), .x(\ILAB0102.ILE0613.net0558 ));
  inv_4_UCCLAB \ILAB0102.ILE0613.I712  ( .a(\ILAB0102.net19976 ), .x(\ILAB0102.ILE0613.net0562 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0714.Ihi5  ( .en(GND), .in(\ILAB0102.ILE0714.net2656 ), .out(\ILAB0102.net19913 ));
  inv_8_UCCLAB \ILAB0102.ILE0716.I666  ( .a(\ILAB0102.net22388 ), .x(\net10355<1> ));
  buf4_12_UCCLAB \ILAB0102.I4397  ( .a(\net10355<1> ), .x(\ILAB0102.net27305 ));
  buftid52C_UCCLAB \ILAB0102.I4458  ( .a(\ILAB0102.net27305 ), .ne(GND), .x(\LongBus_72<14> ));
  buftd52_UCCLAB \ILAB0302.I4801.I26  ( .a(\LongBus_72<14> ), .en(VDD), .x(\LongBus_5<14> ));
  buftd52_UCCLAB \ILAB0303.I4775.I27  ( .a(\LongBus_5<14> ), .en(VDD), .x(\LongBus_71<14> ));
  mux2i_P_UCCLAB \IIO12.I1.I16  ( .d0(GND), .d1(\LongBus_71<14> ), .sl0(VDD), .x(\IIO12.I1.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1204.Ihi5  ( .en(GND), .in(\ILAB0103.ILE1204.net2656 ), .out(\ILAB0103.net26573 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0803.Ivi7  ( .en(GND), .in(\ILAB0103.net26573 ), .out(\ILAB0103.net20344 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0403.Ivi7  ( .en(GND), .in(\ILAB0103.net20344 ), .out(\net11487<6> ));
  inv_8_UCCLAB \ILAB0103.ILE1401.I666  ( .a(\ILAB0103.net26573 ), .x(\net10348<0> ));
  buf4_12_UCCLAB \ILAB0103.I4355  ( .a(\net10348<0> ), .x(\ILAB0103.net39060 ));
  buftid52C_UCCLAB \ILAB0103.I4475  ( .a(\ILAB0103.net39060 ), .ne(GND), .x(\LongBus_71<5> ));
  buftd52_UCCLAB \ILAB0203.I4775.I38  ( .a(\LongBus_71<5> ), .en(VDD), .x(\LongBus_3<5> ));
  buftd52_UCCLAB \ILAB0203.I4801.I39  ( .a(\LongBus_3<5> ), .en(VDD), .x(\LongBus_70<5> ));
  mux2i_P_UCCLAB \IIO12.I2.I16  ( .d0(\LongBus_70<5> ), .d1(GND), .sl0(GND), .x(\IIO12.I2.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1103.Ivi7  ( .en(GND), .in(\ILAB0103.ILE1103.net2656 ), .out(\ILAB0103.net16924 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0703.Ivi7  ( .en(GND), .in(\ILAB0103.net16924 ), .out(\ILAB0103.net15709 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0303.Ivi7  ( .en(GND), .in(\ILAB0103.net15709 ), .out(\net11487<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1103.Ihi5  ( .en(GND), .in(\ILAB0103.ILE1103.net2656 ), .out(\ILAB0103.net16583 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1103.Ivo1  ( .en(GND), .in(\ILAB0103.ILE1103.net2656 ), .out(\ILAB0103.net17734 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1503.Ivo1  ( .en(GND), .in(\ILAB0103.net17734 ), .out(\net18735<3> ));
  inv_8_UCCLAB \ILAB0103.ILE1603.I666  ( .a(\net18735<3> ), .x(\ILAB0103.net26501 ));
  buf4_12_UCCLAB \ILAB0103.I4358  ( .a(\ILAB0103.net26501 ), .x(\ILAB0103.net39588 ));
  buftd52C_UCCLAB \ILAB0103.I4415  ( .a(\ILAB0103.net39588 ), .en(VDD), .x(\LongBus_1<4> ));
  buftd52_UCCLAB \ILAB0103.I4801.I40  ( .a(\LongBus_1<4> ), .en(VDD), .x(\LongBus_70<4> ));
  mux2i_P_UCCLAB \IIO12.I3.I16  ( .d0(\LongBus_70<4> ), .d1(GND), .sl0(GND), .x(\IIO12.I3.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1216.Ihi7  ( .en(GND), .in(\ILAB0102.ILE1216.net2656 ), .out(\ILAB0102.net21352 ));
  inv_8_UCCLAB \ILAB0102.ILE1216.I666  ( .a(\ILAB0102.ILE1216.net0541 ), .x(\net10350<1> ));
  buf4_12_UCCLAB \ILAB0102.I4404  ( .a(\net10350<1> ), .x(\ILAB0102.net27291 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1216.Ivi6  ( .en(GND), .in(\ILAB0102.ILE1216.net2656 ), .out(\ILAB0102.net20974 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0916.Ivi7  ( .en(GND), .in(\ILAB0102.net20974 ), .out(\ILAB0102.net17509 ));
  buftid52C_UCCLAB \ILAB0102.I4461  ( .a(\ILAB0102.net27291 ), .ne(GND), .x(\LongBus_72<11> ));
  buftd52_UCCLAB \ILAB0202.I4801.I22  ( .a(\LongBus_72<11> ), .en(VDD), .x(\LongBus_3<11> ));
  buftd52_UCCLAB \ILAB0203.I4775.I23  ( .a(\LongBus_3<11> ), .en(VDD), .x(\LongBus_71<11> ));
  mux2i_P_UCCLAB \IIO12.I4.I16  ( .d0(GND), .d1(\LongBus_71<11> ), .sl0(VDD), .x(\IIO12.I4.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0813.Ihi7  ( .en(GND), .in(\ILAB0102.ILE0813.net2656 ), .out(\ILAB0102.net17617 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0813.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0813.net2656 ), .out(\ILAB0102.net22549 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0813.Ivo1  ( .en(GND), .in(\ILAB0102.ILE0813.net2656 ), .out(\ILAB0102.net21109 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1213.Ivo1  ( .en(GND), .in(\ILAB0102.net21109 ), .out(\net10337<4> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1613.Ivo1  ( .en(GND), .in(\net10337<4> ), .out(\net18544<6> ));
  inv_8_UCCLAB \ILAB0202.ILE0113.I666  ( .a(\net18544<6> ), .x(\ILAB0202.net21911 ));
  buf4_12_UCCLAB \ILAB0202.I4366  ( .a(\ILAB0202.net21911 ), .x(\ILAB0202.net38625 ));
  buftd52C_UCCLAB \ILAB0202.I4437  ( .a(\ILAB0202.net38625 ), .en(VDD), .x(\LongBus_2<2> ));
  buftd52_UCCLAB \ILAB0203.I4773.I6  ( .a(\LongBus_2<2> ), .en(VDD), .x(\LongBus_70<2> ));
  mux2i_P_UCCLAB \IIO12.I5.I16  ( .d0(\LongBus_70<2> ), .d1(GND), .sl0(GND), .x(\IIO12.I5.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0515.Iho1  ( .en(GND), .in(\ILAB0102.ILE0515.net2656 ), .out(\net10423<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0515.Ivo1  ( .en(GND), .in(\ILAB0102.ILE0515.net2656 ), .out(\ILAB0102.net22189 ));
  inv_8_UCCLAB \ILAB0102.ILE0515.I666  ( .a(\ILAB0102.ILE0515.net0541 ), .x(\ILAB0102.net19796 ));
  inv_4_UCCLAB \ILAB0102.ILE0416.I712  ( .a(\ILAB0102.net19796 ), .x(\ILAB0102.ILE0416.net0562 ));
  inv_4_UCCLAB \ILAB0102.ILE0416.I710  ( .a(\ILAB0102.net19796 ), .x(\ILAB0102.ILE0416.net0558 ));
  inv_8_UCCLAB \ILAB0102.ILE0516.I666  ( .a(\ILAB0102.net19796 ), .x(\net10357<1> ));
  buf4_12_UCCLAB \ILAB0102.I4380  ( .a(\net10357<1> ), .x(\ILAB0102.net27339 ));
  buftid52C_UCCLAB \ILAB0102.I4466  ( .a(\ILAB0102.net27339 ), .ne(GND), .x(\LongBus_72<1> ));
  buftd52_UCCLAB \ILAB0202.I4801.I5  ( .a(\LongBus_72<1> ), .en(VDD), .x(\LongBus_3<1> ));
  buftd52_UCCLAB \ILAB0203.I4801.I4  ( .a(\LongBus_3<1> ), .en(VDD), .x(\LongBus_70<1> ));
  mux2i_P_UCCLAB \IIO12.I6.I16  ( .d0(\LongBus_70<1> ), .d1(GND), .sl0(GND), .x(\IIO12.I6.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1004.Ihi5  ( .en(GND), .in(\ILAB0103.ILE1004.net2656 ), .out(\ILAB0103.net26618 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1004.Ivi7  ( .en(GND), .in(\ILAB0103.ILE1004.net2656 ), .out(\ILAB0103.net23134 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1004.Ivi5  ( .en(GND), .in(\ILAB0103.ILE1004.net2656 ), .out(\ILAB0103.net23132 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1004.Ivo1  ( .en(GND), .in(\ILAB0103.ILE1004.net2656 ), .out(\ILAB0103.net25654 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1404.Ivo1  ( .en(GND), .in(\ILAB0103.net25654 ), .out(\net18731<1> ));
  inv_8_UCCLAB \ILAB0103.ILE1604.I666  ( .a(\net18731<1> ), .x(\ILAB0103.net15476 ));
  buf4_12_UCCLAB \ILAB0103.I4409  ( .a(\ILAB0103.net15476 ), .x(\ILAB0103.net37740 ));
  buftd52C_UCCLAB \ILAB0103.I4430  ( .a(\ILAB0103.net37740 ), .en(VDD), .x(\LongBus_1<0> ));
  buftd52_UCCLAB \ILAB0103.I4801.I1  ( .a(\LongBus_1<0> ), .en(VDD), .x(\LongBus_70<0> ));
  mux2i_P_UCCLAB \IIO12.I7.I16  ( .d0(\LongBus_70<0> ), .d1(GND), .sl0(GND), .x(\IIO12.I7.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0602.Ivo1  ( .en(GND), .in(\ILAB0103.ILE0602.net2656 ), .out(\ILAB0103.net26644 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0602.Ihi5  ( .en(GND), .in(\ILAB0103.ILE0602.net2656 ), .out(\net10419<5> ));
  inv_8_UCCLAB \ILAB0103.ILE0602.I666  ( .a(\ILAB0103.ILE0602.net0541 ), .x(\ILAB0103.net20606 ));
  inv_4_UCCLAB \ILAB0103.ILE0701.I714  ( .a(\ILAB0103.net20606 ), .x(\ILAB0103.ILE0701.net01345 ));
  inv_8_UCCLAB \ILAB0103.ILE0601.I666  ( .a(\ILAB0103.net20606 ), .x(\net10356<0> ));
  buf4_12_UCCLAB \ILAB0103.I4412  ( .a(\net10356<0> ), .x(\ILAB0103.net38382 ));
  buftid52C_UCCLAB \ILAB0103.I4476  ( .a(\ILAB0103.net38382 ), .ne(GND), .x(\LongBus_71<15> ));
  buftd52_UCCLAB \ILAB0203.I4772.I29  ( .a(\LongBus_71<15> ), .en(VDD), .x(\LongBus_2<15> ));
  buftd52_UCCLAB \ILAB0204.I4772.I28  ( .a(\LongBus_2<15> ), .en(VDD), .x(\LongBus_69<15> ));
  mux2i_P_UCCLAB \IIO13.I0.I16  ( .d0(GND), .d1(\LongBus_69<15> ), .sl0(VDD), .x(\IIO13.I0.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0503.Ihi5  ( .en(GND), .in(\ILAB0103.ILE0503.net2656 ), .out(\ILAB0103.net20633 ));
  inv_8_UCCLAB \ILAB0103.ILE0503.I666  ( .a(\ILAB0103.ILE0503.net0541 ), .x(\ILAB0103.net26276 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0503.Ivi5  ( .en(GND), .in(\ILAB0103.ILE0503.net2656 ), .out(\ILAB0103.net20162 ));
  inv_4_UCCLAB \ILAB0103.ILE0402.I710  ( .a(\ILAB0103.net26276 ), .x(\ILAB0103.ILE0402.net0558 ));
  inv_4_UCCLAB \ILAB0103.ILE0402.I712  ( .a(\ILAB0103.net26276 ), .x(\ILAB0103.ILE0402.net0562 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0503.Ivi7  ( .en(GND), .in(\ILAB0103.ILE0503.net2656 ), .out(\Fast_out_29<5> ));
  inv_8_UCCLAB \ILAB0103.ILE0105.I666  ( .a(\Fast_out_29<5> ), .x(\ILAB0103.net22946 ));
  buf4_12_UCCLAB \ILAB0103.I4379  ( .a(\ILAB0103.net22946 ), .x(\ILAB0103.net38496 ));
  buftd52C_UCCLAB \ILAB0103.I4441  ( .a(\ILAB0103.net38496 ), .en(VDD), .x(\LongBus_0<14> ));
  buftd52_UCCLAB \ILAB0104.I4772.I27  ( .a(\LongBus_0<14> ), .en(VDD), .x(\LongBus_69<14> ));
  mux2i_P_UCCLAB \IIO13.I1.I16  ( .d0(GND), .d1(\LongBus_69<14> ), .sl0(VDD), .x(\IIO13.I1.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0904.Ihi5  ( .en(GND), .in(\ILAB0103.ILE0904.net2656 ), .out(\ILAB0103.net26168 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0904.Ivi7  ( .en(GND), .in(\ILAB0103.ILE0904.net2656 ), .out(\ILAB0103.net25114 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0904.Ivi5  ( .en(GND), .in(\ILAB0103.ILE0904.net2656 ), .out(\ILAB0103.net25112 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0704.Ivi6  ( .en(GND), .in(\ILAB0103.net25112 ), .out(\ILAB0103.net25609 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0404.Ivi7  ( .en(GND), .in(\ILAB0103.net25609 ), .out(\net11483<6> ));
  inv_8_UCCLAB \ILAB0103.ILE0104.I666  ( .a(\net11483<6> ), .x(\ILAB0103.net22856 ));
  buf4_12_UCCLAB \ILAB0103.I4378  ( .a(\ILAB0103.net22856 ), .x(\ILAB0103.net37425 ));
  buftd52C_UCCLAB \ILAB0103.I4434  ( .a(\ILAB0103.net37425 ), .en(VDD), .x(\LongBus_0<5> ));
  buftd52_UCCLAB \ILAB0104.I4773.I39  ( .a(\LongBus_0<5> ), .en(VDD), .x(\LongBus_68<5> ));
  mux2i_P_UCCLAB \IIO13.I2.I16  ( .d0(\LongBus_68<5> ), .d1(GND), .sl0(GND), .x(\IIO13.I2.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0704.Ihi5  ( .en(GND), .in(\ILAB0103.ILE0704.net2656 ), .out(\ILAB0103.net26438 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0704.Ihi7  ( .en(GND), .in(\ILAB0103.ILE0704.net2656 ), .out(\net10415<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0704.Ivi7  ( .en(GND), .in(\ILAB0103.ILE0704.net2656 ), .out(\ILAB0103.net16114 ));
  inv_8_UCCLAB \ILAB0103.ILE0701.I666  ( .a(\net10415<6> ), .x(\net10355<0> ));
  buf4_12_UCCLAB \ILAB0103.I4395  ( .a(\net10355<0> ), .x(\ILAB0103.net39618 ));
  buftid52C_UCCLAB \ILAB0103.I4473  ( .a(\ILAB0103.net39618 ), .ne(GND), .x(\LongBus_71<4> ));
  buftd52_UCCLAB \ILAB0203.I4775.I41  ( .a(\LongBus_71<4> ), .en(VDD), .x(\LongBus_3<4> ));
  buftd52_UCCLAB \ILAB0204.I4801.I40  ( .a(\LongBus_3<4> ), .en(VDD), .x(\LongBus_68<4> ));
  mux2i_P_UCCLAB \IIO13.I3.I16  ( .d0(\LongBus_68<4> ), .d1(GND), .sl0(GND), .x(\IIO13.I3.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0401.Ivi7  ( .en(GND), .in(\ILAB0103.ILE0401.net2656 ), .out(\net11495<6> ));
  inv_8_UCCLAB \ILAB0103.ILE0401.I666  ( .a(\ILAB0103.ILE0401.net0541 ), .x(\net10358<0> ));
  buf4_12_UCCLAB \ILAB0103.I4411  ( .a(\net10358<0> ), .x(\ILAB0103.net37923 ));
  buftid52C_UCCLAB \ILAB0103.I4474  ( .a(\ILAB0103.net37923 ), .ne(GND), .x(\LongBus_71<3> ));
  buftd52_UCCLAB \ILAB0203.I4772.I9  ( .a(\LongBus_71<3> ), .en(VDD), .x(\LongBus_2<3> ));
  buftd52_UCCLAB \ILAB0204.I4773.I8  ( .a(\LongBus_2<3> ), .en(VDD), .x(\LongBus_68<3> ));
  mux2i_P_UCCLAB \IIO13.I4.I16  ( .d0(\LongBus_68<3> ), .d1(GND), .sl0(GND), .x(\IIO13.I4.net197 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0401.Ivo2  ( .en(GND), .in(\ILAB0103.ILE0401.net2656 ), .out(\ILAB0103.net20612 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0611.Ivo1  ( .en(GND), .in(\ILAB0102.ILE0611.net2656 ), .out(\ILAB0102.net22684 ));
  inv_8_UCCLAB \ILAB0102.ILE0611.I666  ( .a(\ILAB0102.ILE0611.net0541 ), .x(\ILAB0102.net24116 ));
  inv_4_UCCLAB \ILAB0102.ILE0510.I712  ( .a(\ILAB0102.net24116 ), .x(\ILAB0102.ILE0510.net0562 ));
  inv_4_UCCLAB \ILAB0102.ILE0510.I710  ( .a(\ILAB0102.net24116 ), .x(\ILAB0102.ILE0510.net0558 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0611.Ivi5  ( .en(GND), .in(\ILAB0102.ILE0611.net2656 ), .out(\ILAB0102.net21467 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1011.Ivo1  ( .en(GND), .in(\ILAB0102.net22684 ), .out(\ILAB0102.net20434 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1411.Ivo1  ( .en(GND), .in(\ILAB0102.net20434 ), .out(\net18552<1> ));
  inv_8_UCCLAB \ILAB0102.ILE1611.I666  ( .a(\net18552<1> ), .x(\ILAB0102.net24386 ));
  buf4_12_UCCLAB \ILAB0102.I4399  ( .a(\ILAB0102.net24386 ), .x(\ILAB0102.net38760 ));
  buftd52C_UCCLAB \ILAB0102.I4422  ( .a(\ILAB0102.net38760 ), .en(VDD), .x(\LongBus_1<2> ));
  buftd52_UCCLAB \ILAB0104.I4801.I6  ( .a(\LongBus_1<2> ), .en(VDD), .x(\LongBus_68<2> ));
  mux2i_P_UCCLAB \IIO13.I5.I16  ( .d0(\LongBus_68<2> ), .d1(GND), .sl0(GND), .x(\IIO13.I5.net197 ));
  mux4p_0_UCCLAB \IIO31.I24  ( .d0(\Fast_in_32<7> ), .d1(GND), .d2(GND), .d3(GND), .sl0(GND), .sl1(GND), .x(\IIO31.net728 ));
  invtd56_clk1_UCCLAB \IIO31.I12  ( .a(\IIO31.net728 ), .en(VDD), .x(\net9202<2> ));
  mux4p_0_AVDD \I3621.I152.I13  ( .d0(GND), .d1(GND), .d2(GND), .d3(\net9202<2> ), .sl0(VDD), .sl1(VDD), .x(\I3621.I152.net117 ));
  invtd56_pd_clk_AVDD \I3621.I152.I5  ( .a(\I3621.I152.net117 ), .en(VDD), .x(\net10329<2> ));
  mux4p_0_UCCLAB \I3590.I13  ( .d0(GND), .d1(\net10329<2> ), .d2(GND), .d3(GND), .sl0(VDD), .sl1(GND), .x(\I3590.net78 ));
  invtd56_pd_clk_UCCLAB \I3590.I5  ( .a(\I3590.net78 ), .en(VDD), .x(\net10262<1> ));
  mux2p_2_UCCLAB \I3687.I4  ( .d0(\net10262<1> ), .d1(GND), .s0(GND), .x(\I3687.net43 ));
  invtd56_pd_clk_UCCLAB \I3687.I5  ( .a(\I3687.net43 ), .en(VDD), .x(\net21016<1> ));
  invtd56_pd_clk_UCCLAB \I3635.I2  ( .a(\net21016<1> ), .en(VDD), .x(\GCLK_s5<2> ));
  nand2_1_UCCLAB \ILAB1001.I5366.I72  ( .a(VDD), .b(\GCLK_s5<2> ), .x(\ILAB1001.I5366.net68 ));
  mux2d1i_1_P_UCCLAB \ILAB1001.I5366.I80  ( .d0(GND), .d1i(\ILAB1001.I5366.net68 ), .sl0(VDD), .x(\ILAB1001.I5366.net0106 ));
  invd52_UCCLAB \ILAB1001.I5366.I76  ( .a(\ILAB1001.I5366.net0106 ), .x(\ILAB1001.net15299<1> ));
  invd32_UCCLAB \ILAB1001.I5591.I1  ( .a(\ILAB1001.net15299<1> ), .x(\ILAB1001.Clk_LAB<2> ));
  sw_b_v2_inv_UCCLAB \ILAB1001.ILE1403.Iho1  ( .en(GND), .in(\ILAB1001.ILE1403.net2656 ), .out(\ILAB1001.net20002 ));
  sw_b_v2_inv_UCCLAB \ILAB1001.ILE1407.Iho1  ( .en(GND), .in(\ILAB1001.net20002 ), .out(\ILAB1001.net25762 ));
  sw_b_v2_inv_UCCLAB \ILAB0201.ILE0314.Ihi7  ( .en(GND), .in(\ILAB0201.ILE0314.net2656 ), .out(\ILAB0201.net25897 ));
  sw_b_v2_inv_UCCLAB \ILAB0201.ILE0314.Ivi6  ( .en(GND), .in(\ILAB0201.ILE0314.net2656 ), .out(\net18389<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0201.ILE0314.Ivi5  ( .en(GND), .in(\ILAB0201.ILE0314.net2656 ), .out(\ILAB0201.net23807 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1602.Iho1  ( .en(GND), .in(\net18389<6> ), .out(\ILAB0102.net26482 ));
  sw_b_v2_inv_UCCLAB \ILAB0101.ILE1613.Ivi7  ( .en(GND), .in(\ILAB0201.net25897 ), .out(\net17132<4> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1605.Iho2  ( .en(GND), .in(\ILAB0102.net26482 ), .out(\ILAB0102.net15863 ));
  sw_b_v2_inv_UCCLAB \ILAB0202.ILE0101.Iho2  ( .en(GND), .in(\ILAB0201.net23807 ), .out(\ILAB0202.net16718 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1405.Ivi6  ( .en(GND), .in(\ILAB0102.net26482 ), .out(\ILAB0102.net15754 ));
  sw_b_v2_inv_UCCLAB \ILAB0202.ILE0205.Ivi6  ( .en(GND), .in(\ILAB0202.ILE0205.net2656 ), .out(\net18576<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0101.ILE1513.Iho1  ( .en(GND), .in(\ILAB0101.ILE1513.net2656 ), .out(\net17178<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1501.Iho1  ( .en(GND), .in(\net17178<0> ), .out(\ILAB0102.net20857 ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0202.Ivo1  ( .en(GND), .in(\ILAB0402.ILE0202.net2656 ), .out(\ILAB0402.net26419 ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0202.Ihi5  ( .en(GND), .in(\ILAB0402.ILE0202.net2656 ), .out(\net16324<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0202.Ihi7  ( .en(GND), .in(\ILAB0402.ILE0202.net2656 ), .out(\net16324<1> ));
  inv_8_UCCLAB \ILAB0402.ILE0202.I666  ( .a(\ILAB0402.ILE0202.net0541 ), .x(\ILAB0402.net16961 ));
  inv_4_UCCLAB \ILAB0402.ILE0301.I715  ( .a(\ILAB0402.net16961 ), .x(\ILAB0402.ILE0301.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0313.Iho3  ( .en(GND), .in(\ILAB0401.ILE0313.net2656 ), .out(\ILAB0401.net23154 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0313.Iho2  ( .en(GND), .in(\ILAB0401.ILE0313.net2656 ), .out(\ILAB0401.net23153 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0313.Ivi5  ( .en(GND), .in(\ILAB0401.ILE0313.net2656 ), .out(\ILAB0401.net23177 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0313.Ivi7  ( .en(GND), .in(\ILAB0401.ILE0313.net2656 ), .out(\net16279<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0213.Ivo2  ( .en(GND), .in(\net16279<3> ), .out(\ILAB0401.net26102 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0314.Ivo1  ( .en(GND), .in(\ILAB0401.ILE0314.net2656 ), .out(\ILAB0401.net22414 ));
  inv_8_UCCLAB \ILAB0401.ILE0514.I666  ( .a(\ILAB0401.net22414 ), .x(\ILAB0401.net18311 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0113.Iho2  ( .en(GND), .in(\ILAB0401.ILE0113.net2656 ), .out(\ILAB0401.net22253 ));
  inv_8_UCCLAB \ILAB0401.ILE0113.I666  ( .a(\ILAB0401.ILE0113.net0541 ), .x(\ILAB0401.net21911 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0115.Iho3  ( .en(GND), .in(\ILAB0401.net22253 ), .out(\ILAB0401.net24549 ));
  inv_4_UCCLAB \ILAB0401.ILE0214.I715  ( .a(\ILAB0401.net21911 ), .x(\ILAB0401.ILE0214.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0113.Iho3  ( .en(GND), .in(\ILAB0401.ILE0113.net2656 ), .out(\ILAB0401.net22254 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0113.Ivo1  ( .en(GND), .in(\ILAB0401.ILE0113.net2656 ), .out(\ILAB0401.net18319 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0214.Ivo1  ( .en(GND), .in(\ILAB0401.net22254 ), .out(\ILAB0401.net22144 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0312.Iho1  ( .en(GND), .in(\ILAB0401.ILE0312.net2656 ), .out(\ILAB0401.net24907 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0312.Ivo1  ( .en(GND), .in(\ILAB0401.ILE0312.net2656 ), .out(\ILAB0401.net19939 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0312.Ivi7  ( .en(GND), .in(\ILAB0401.ILE0312.net2656 ), .out(\net16283<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0312.Iho2  ( .en(GND), .in(\ILAB0401.ILE0312.net2656 ), .out(\ILAB0401.net24908 ));
  inv_8_UCCLAB \ILAB0401.ILE0312.I666  ( .a(\ILAB0401.ILE0312.net0541 ), .x(\ILAB0401.net23396 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0314.Iho3  ( .en(GND), .in(\ILAB0401.net24908 ), .out(\ILAB0401.net23784 ));
  inv_4_UCCLAB \ILAB0401.ILE0413.I714  ( .a(\ILAB0401.net23396 ), .x(\ILAB0401.ILE0413.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0413.Ivo3  ( .en(GND), .in(\ILAB0401.ILE0413.net2656 ), .out(\ILAB0401.net18315 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0215.Ivi7  ( .en(GND), .in(\ILAB0401.ILE0215.net2656 ), .out(\net16271<1> ));
  inv_8_UCCLAB \ILAB0301.ILE1615.I666  ( .a(\net16271<1> ), .x(\ILAB0301.net22766 ));
  buftd4_UCCLAB \ILAB0301.I180  ( .a(\ILAB0301.net22766 ), .en(VDD), .x(\ILAB0301.net015234 ));
  mux2p_2_UCCLAB \ILAB0301.I5605.I0  ( .d0(GND), .d1(\ILAB0301.net015234 ), .s0(VDD), .x(\ILAB0301.I5605.net29 ));
  invd16_seth_UCCLAB \ILAB0301.I5605.I1  ( .a(\ILAB0301.I5605.net29 ), .c(VDD), .x(\ILAB0301.Clk_int<3> ));
  mux2p_2_UCCLAB \ILAB0301.I5366.I83  ( .d0(GND), .d1(\ILAB0301.Clk_int<3> ), .s0(VDD), .x(\ILAB0301.I5366.net0122 ));
  invtd56_clk_UCCLAB \ILAB0301.I5366.I8  ( .a(\ILAB0301.I5366.net0122 ), .en(VDD), .x(\net16372<0> ));
  invtd56_UCCLAB \I3700.I3  ( .a(\net16372<0> ), .en(VDD), .x(\net10281<0> ));
  mux2p_2_UCCLAB \I3690.I3  ( .d0(GND), .d1(\net10281<0> ), .s0(VDD), .x(\I3690.net39 ));
  invtd56_pd_clk_UCCLAB \I3690.I7  ( .a(\I3690.net39 ), .en(VDD), .x(\net20974<2> ));
  invtd56_pd_clk_UCCLAB \I3651.I3  ( .a(\net20974<2> ), .en(VDD), .x(\GCLK_s1<1> ));
  nand2_1_UCCLAB \ILAB0202.I5366.I71  ( .a(VDD), .b(\GCLK_s1<1> ), .x(\ILAB0202.I5366.net70 ));
  mux2d1i_1_P_UCCLAB \ILAB0202.I5366.I79  ( .d0(GND), .d1i(\ILAB0202.I5366.net70 ), .sl0(VDD), .x(\ILAB0202.I5366.net0110 ));
  invd52_UCCLAB \ILAB0202.I5366.I75  ( .a(\ILAB0202.I5366.net0110 ), .x(\ILAB0202.net15299<2> ));
  invd32_UCCLAB \ILAB0202.I5591.I2  ( .a(\ILAB0202.net15299<2> ), .x(\ILAB0202.Clk_LAB<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0502.Ihi5  ( .en(GND), .in(\ILAB0402.ILE0502.net2656 ), .out(\net16312<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0502.Ivi7  ( .en(GND), .in(\ILAB0402.ILE0502.net2656 ), .out(\net11247<1> ));
  inv_8_UCCLAB \ILAB0402.ILE0502.I666  ( .a(\ILAB0402.ILE0502.net0541 ), .x(\ILAB0402.net20651 ));
  inv_4_UCCLAB \ILAB0402.ILE0401.I712  ( .a(\ILAB0402.net20651 ), .x(\ILAB0402.ILE0401.net0562 ));
  inv_4_UCCLAB \ILAB0402.ILE0401.I710  ( .a(\ILAB0402.net20651 ), .x(\ILAB0402.ILE0401.net0558 ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0502.Ihi6  ( .en(GND), .in(\ILAB0402.ILE0502.net2656 ), .out(\net16312<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0716.Ivi7  ( .en(GND), .in(\ILAB0401.ILE0716.net2656 ), .out(\ILAB0401.net19309 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0716.Iho2  ( .en(GND), .in(\ILAB0401.ILE0716.net2656 ), .out(\net16304<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0302.Ivi6  ( .en(GND), .in(\ILAB0402.ILE0302.net2656 ), .out(\net11340<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0302.ILE1602.Ivi7  ( .en(GND), .in(\net11340<6> ), .out(\ILAB0302.net26509 ));
  sw_b_v2_inv_UCCLAB \ILAB0302.ILE1202.Ivi7  ( .en(GND), .in(\ILAB0302.net26509 ), .out(\ILAB0302.net26599 ));
  sw_b_v2_inv_UCCLAB \ILAB0302.ILE0802.Ivi7  ( .en(GND), .in(\ILAB0302.net26599 ), .out(\ILAB0302.net26149 ));
  sw_b_v2_inv_UCCLAB \ILAB0302.ILE0402.Ivi7  ( .en(GND), .in(\ILAB0302.net26149 ), .out(\net11189<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0202.ILE1602.Ivi7  ( .en(GND), .in(\net11189<6> ), .out(\ILAB0202.net26509 ));
  sw_b_v2_inv_UCCLAB \ILAB0202.ILE1202.Ivi7  ( .en(GND), .in(\ILAB0202.net26509 ), .out(\ILAB0202.net26599 ));
  sw_b_v2_inv_UCCLAB \ILAB0202.ILE0802.Ivi7  ( .en(GND), .in(\ILAB0202.net26599 ), .out(\ILAB0202.net26149 ));
  sw_b_v2_inv_UCCLAB \ILAB0202.ILE0402.Ivi7  ( .en(GND), .in(\ILAB0202.net26149 ), .out(\net18588<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0202.ILE0202.Ivi7  ( .en(GND), .in(\ILAB0202.ILE0202.net2656 ), .out(\net18588<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0202.ILE0202.Ivi5  ( .en(GND), .in(\ILAB0202.ILE0202.net2656 ), .out(\net18588<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1602.Ivi6  ( .en(GND), .in(\net18588<5> ), .out(\net18588<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1302.Ivi7  ( .en(GND), .in(\net18588<0> ), .out(\ILAB0102.net26554 ));
  sw_b_v2_inv_UCCLAB \ILAB0302.ILE1501.Ivo1  ( .en(GND), .in(\ILAB0302.ILE1501.net2656 ), .out(\net11344<3> ));
  inv_8_UCCLAB \ILAB0302.ILE1501.I666  ( .a(\ILAB0302.ILE1501.net0541 ), .x(\net16387<0> ));
  buf4_12_UCCLAB \ILAB0302.I4368  ( .a(\net16387<0> ), .x(\ILAB0302.net38580 ));
  buftid52C_UCCLAB \ILAB0302.I4477  ( .a(\ILAB0302.net38580 ), .ne(GND), .x(\LongBus_73<0> ));
  buftid52C_UCCLAB \ILAB0302.I4457  ( .a(\ILAB0302.net38580 ), .ne(GND), .x(\LongBus_73<1> ));
  buftd52_UCCLAB \ILAB0102.I4775.I5  ( .a(\LongBus_73<1> ), .en(VDD), .x(\LongBus_1<1> ));
  buftd52_UCCLAB \ILAB0202.I4772.I62895  ( .a(\LongBus_73<0> ), .en(VDD), .x(\LongBus_2<0> ));
  inv_8_UCCLAB \ILAB0302.ILE1601.I666  ( .a(\net11344<3> ), .x(\net16386<0> ));
  buftd4_UCCLAB \ILAB0302.I237  ( .a(\net16386<0> ), .en(VDD), .x(\ILAB0302.net027160 ));
  mux2p_2_UCCLAB \ILAB0302.I5605.I7  ( .d0(\ILAB0302.net027160 ), .d1(GND), .s0(GND), .x(\ILAB0302.I5605.net21 ));
  invd16_seth_UCCLAB \ILAB0302.I5605.I6  ( .a(\ILAB0302.I5605.net21 ), .c(VDD), .x(\ILAB0302.Clk_int<0> ));
  mux2p_2_UCCLAB \ILAB0302.I5366.I82  ( .d0(\ILAB0302.Clk_int<0> ), .d1(GND), .s0(GND), .x(\ILAB0302.I5366.net0119 ));
  invtd56_clk_UCCLAB \ILAB0302.I5366.I6  ( .a(\ILAB0302.I5366.net0119 ), .en(VDD), .x(\net16372<1> ));
  inv_4_UCCLAB \ILAB0102.ILE1604.I710  ( .a(\LongBus_1<1> ), .x(\ILAB0102.ILE1604.net0558 ));
  inv_4_UCCLAB \ILAB0202.ILE0103.I713  ( .a(\LongBus_2<0> ), .x(\ILAB0202.ILE0103.net01342 ));
  invtd56_UCCLAB \I3700.I4  ( .a(\net16372<1> ), .en(VDD), .x(\net10281<1> ));
  mux2p_2_UCCLAB \I3690.I4  ( .d0(GND), .d1(\net10281<1> ), .s0(VDD), .x(\I3690.net43 ));
  invtd56_pd_clk_UCCLAB \I3690.I5  ( .a(\I3690.net43 ), .en(VDD), .x(\net20974<1> ));
  invtd56_pd_clk_UCCLAB \I3651.I2  ( .a(\net20974<1> ), .en(VDD), .x(\GCLK_s1<2> ));
  nand2_1_UCCLAB \ILAB0202.I5366.I72  ( .a(VDD), .b(\GCLK_s1<2> ), .x(\ILAB0202.I5366.net68 ));
  mux2d1i_1_P_UCCLAB \ILAB0202.I5366.I80  ( .d0(GND), .d1i(\ILAB0202.I5366.net68 ), .sl0(VDD), .x(\ILAB0202.I5366.net0106 ));
  invd52_UCCLAB \ILAB0202.I5366.I76  ( .a(\ILAB0202.I5366.net0106 ), .x(\ILAB0202.net15299<1> ));
  invd32_UCCLAB \ILAB0202.I5591.I1  ( .a(\ILAB0202.net15299<1> ), .x(\ILAB0202.Clk_LAB<2> ));
  nand2_1_UCCLAB \ILAB0102.I5366.I72  ( .a(VDD), .b(\GCLK_s1<2> ), .x(\ILAB0102.I5366.net68 ));
  mux2d1i_1_P_UCCLAB \ILAB0102.I5366.I80  ( .d0(GND), .d1i(\ILAB0102.I5366.net68 ), .sl0(VDD), .x(\ILAB0102.I5366.net0106 ));
  invd52_UCCLAB \ILAB0102.I5366.I76  ( .a(\ILAB0102.I5366.net0106 ), .x(\ILAB0102.net15299<1> ));
  invd32_UCCLAB \ILAB0102.I5591.I1  ( .a(\ILAB0102.net15299<1> ), .x(\ILAB0102.Clk_LAB<2> ));
  sw_b_v2_inv_UCCLAB \ILAB0202.ILE0302.Ivi7  ( .en(GND), .in(\ILAB0202.ILE0302.net2656 ), .out(\net18588<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0202.ILE0302.Ivi5  ( .en(GND), .in(\ILAB0202.ILE0302.net2656 ), .out(\ILAB0202.net26822 ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0102.Ihi7  ( .en(GND), .in(\ILAB0402.ILE0102.net2656 ), .out(\net16328<1> ));
  inv_8_UCCLAB \ILAB0402.ILE0102.I666  ( .a(\ILAB0402.ILE0102.net0541 ), .x(\ILAB0402.net16736 ));
  buf4_12_UCCLAB \ILAB0402.I4388  ( .a(\ILAB0402.net16736 ), .x(\ILAB0402.net37806 ));
  buftd52C_UCCLAB \ILAB0402.I4443  ( .a(\ILAB0402.net37806 ), .en(VDD), .x(\LongBus_6<4> ));
  buftd52_UCCLAB \ILAB0402.I4772.I40  ( .a(\LongBus_6<4> ), .en(VDD), .x(\net8296<11> ));
  buftd52C_UCCLAB \I3741.I41  ( .a(\net8296<11> ), .en(VDD), .x(\LongBus_73<4> ));
  buftd52_UCCLAB \ILAB0202.I4772.I41  ( .a(\LongBus_73<4> ), .en(VDD), .x(\LongBus_2<4> ));
  inv_4_UCCLAB \ILAB0202.ILE0103.I714  ( .a(\LongBus_2<4> ), .x(\ILAB0202.ILE0103.net01345 ));
  buftd52C_UCCLAB \ILAB0402.I4434  ( .a(\ILAB0402.net37806 ), .en(VDD), .x(\LongBus_6<5> ));
  buftd52_UCCLAB \ILAB0402.I4772.I39  ( .a(\LongBus_6<5> ), .en(VDD), .x(\net8296<10> ));
  buftd52C_UCCLAB \I3741.I38  ( .a(\net8296<10> ), .en(VDD), .x(\LongBus_73<5> ));
  inv_4_UCCLAB \ILAB0102.ILE1401.I715  ( .a(\LongBus_73<5> ), .x(\ILAB0102.ILE1401.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1402.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1402.net2656 ), .out(\ILAB0102.net26329 ));
  inv_8_UCCLAB \ILAB0102.ILE1402.I666  ( .a(\ILAB0102.ILE1402.net0541 ), .x(\ILAB0102.net20831 ));
  inv_4_UCCLAB \ILAB0102.ILE1303.I711  ( .a(\ILAB0102.net20831 ), .x(\ILAB0102.ILE1303.net0560 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1403.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1403.net2656 ), .out(\ILAB0102.net20029 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1403.Ivo2  ( .en(GND), .in(\ILAB0102.ILE1403.net2656 ), .out(\ILAB0102.net15482 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1403.Ihi6  ( .en(GND), .in(\ILAB0102.ILE1403.net2656 ), .out(\net17182<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1404.Iho1  ( .en(GND), .in(\net17182<6> ), .out(\ILAB0102.net25627 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1408.Iho1  ( .en(GND), .in(\ILAB0102.net25627 ), .out(\ILAB0102.net19507 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1005.Iho3  ( .en(GND), .in(\ILAB0102.net20029 ), .out(\ILAB0102.net17799 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1412.Iho1  ( .en(GND), .in(\ILAB0102.net19507 ), .out(\ILAB0102.net19372 ));
  inv_8_UCCLAB \ILAB0102.ILE1603.I666  ( .a(\ILAB0102.net15482 ), .x(\ILAB0102.net26501 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1503.Iho1  ( .en(GND), .in(\ILAB0102.net15482 ), .out(\ILAB0102.net17707 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1007.Iho1  ( .en(GND), .in(\ILAB0102.net20029 ), .out(\ILAB0102.net25807 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1507.Iho1  ( .en(GND), .in(\ILAB0102.net17707 ), .out(\ILAB0102.net25717 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1011.Iho1  ( .en(GND), .in(\ILAB0102.net25807 ), .out(\ILAB0102.net22657 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0905.Ivo2  ( .en(GND), .in(\ILAB0102.net20029 ), .out(\ILAB0102.net17957 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1416.Iho1  ( .en(GND), .in(\ILAB0102.net19372 ), .out(\net10387<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1511.Iho1  ( .en(GND), .in(\ILAB0102.net25717 ), .out(\ILAB0102.net21262 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1015.Iho1  ( .en(GND), .in(\ILAB0102.net22657 ), .out(\net10403<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1514.Iho2  ( .en(GND), .in(\ILAB0102.net21262 ), .out(\ILAB0102.net22028 ));
  buftd4_UCCLAB \ILAB0102.I227  ( .a(\ILAB0102.net26501 ), .en(VDD), .x(\ILAB0102.net027166 ));
  mux2p_2_UCCLAB \ILAB0102.I5605.I4  ( .d0(\ILAB0102.net027166 ), .d1(GND), .s0(GND), .x(\ILAB0102.I5605.net25 ));
  invd16_seth_UCCLAB \ILAB0102.I5605.I5  ( .a(\ILAB0102.I5605.net25 ), .c(VDD), .x(\ILAB0102.Clk_int<1> ));
  mux2d1i_1_P_UCCLAB \ILAB0102.I5366.I79  ( .d0(\ILAB0102.Clk_int<1> ), .d1i(GND), .sl0(GND), .x(\ILAB0102.I5366.net0110 ));
  invd52_UCCLAB \ILAB0102.I5366.I75  ( .a(\ILAB0102.I5366.net0110 ), .x(\ILAB0102.net15299<2> ));
  invd32_UCCLAB \ILAB0102.I5591.I2  ( .a(\ILAB0102.net15299<2> ), .x(\ILAB0102.Clk_LAB<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0202.ILE0103.Iho1  ( .en(GND), .in(\ILAB0202.ILE0103.net2656 ), .out(\ILAB0202.net22837 ));
  sw_b_v2_inv_UCCLAB \ILAB0202.ILE0103.Ivi6  ( .en(GND), .in(\ILAB0202.ILE0103.net2656 ), .out(\net18584<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0202.ILE0103.Ivi5  ( .en(GND), .in(\ILAB0202.ILE0103.net2656 ), .out(\net18584<2> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1502.Iho3  ( .en(GND), .in(\ILAB0102.ILE1502.net2656 ), .out(\ILAB0102.net26349 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1103.Ivi7  ( .en(GND), .in(\ILAB0102.net26349 ), .out(\ILAB0102.net16924 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0703.Ivi7  ( .en(GND), .in(\ILAB0102.net16924 ), .out(\ILAB0102.net15709 ));
  inv_8_UCCLAB \ILAB0102.ILE1503.I666  ( .a(\ILAB0102.ILE1503.net0541 ), .x(\ILAB0102.net26366 ));
  inv_4_UCCLAB \ILAB0102.ILE1602.I715  ( .a(\ILAB0102.net26366 ), .x(\ILAB0102.ILE1602.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1602.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1602.net2656 ), .out(\ILAB0102.net26509 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1303.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1303.net2656 ), .out(\ILAB0102.net16654 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1303.Ivi5  ( .en(GND), .in(\ILAB0102.ILE1303.net2656 ), .out(\ILAB0102.net16652 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1303.Iho1  ( .en(GND), .in(\ILAB0102.ILE1303.net2656 ), .out(\ILAB0102.net16627 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0906.Iho2  ( .en(GND), .in(\ILAB0102.net16654 ), .out(\ILAB0102.net24638 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1107.Iho1  ( .en(GND), .in(\ILAB0102.net16652 ), .out(\ILAB0102.net17167 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1001.Ihi6  ( .en(GND), .in(\ILAB0102.net16654 ), .out(\net17198<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1307.Iho1  ( .en(GND), .in(\ILAB0102.net16627 ), .out(\ILAB0102.net17122 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1002.Iho1  ( .en(GND), .in(\net17198<1> ), .out(\ILAB0102.net26617 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1111.Iho1  ( .en(GND), .in(\ILAB0102.net17167 ), .out(\ILAB0102.net23017 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1311.Iho1  ( .en(GND), .in(\ILAB0102.net17122 ), .out(\ILAB0102.net22207 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1006.Iho1  ( .en(GND), .in(\ILAB0102.net26617 ), .out(\ILAB0102.net18202 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1115.Iho1  ( .en(GND), .in(\ILAB0102.net23017 ), .out(\net10399<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1314.Iho2  ( .en(GND), .in(\ILAB0102.net22207 ), .out(\ILAB0102.net23243 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0909.Iho1  ( .en(GND), .in(\ILAB0102.net24638 ), .out(\ILAB0102.net25312 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0913.Iho1  ( .en(GND), .in(\ILAB0102.net25312 ), .out(\net10407<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1010.Iho1  ( .en(GND), .in(\ILAB0102.net18202 ), .out(\ILAB0102.net24862 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1014.Iho1  ( .en(GND), .in(\ILAB0102.net24862 ), .out(\net10403<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1304.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1304.net2656 ), .out(\ILAB0102.net25159 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1304.Iho2  ( .en(GND), .in(\ILAB0102.ILE1304.net2656 ), .out(\ILAB0102.net25133 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0904.Ivi7  ( .en(GND), .in(\ILAB0102.net25159 ), .out(\ILAB0102.net25114 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0908.Iho1  ( .en(GND), .in(\ILAB0102.net25159 ), .out(\ILAB0102.net18517 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1105.Iho1  ( .en(GND), .in(\ILAB0102.net25159 ), .out(\ILAB0102.net17932 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1109.Iho1  ( .en(GND), .in(\ILAB0102.net17932 ), .out(\ILAB0102.net16357 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1113.Iho1  ( .en(GND), .in(\ILAB0102.net16357 ), .out(\net10399<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1304.Ihi6  ( .en(GND), .in(\ILAB0102.ILE1304.net2656 ), .out(\ILAB0102.net20452 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1305.Iho1  ( .en(GND), .in(\ILAB0102.net20452 ), .out(\ILAB0102.net15907 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1309.Iho1  ( .en(GND), .in(\ILAB0102.net15907 ), .out(\ILAB0102.net16222 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1313.Iho1  ( .en(GND), .in(\ILAB0102.net16222 ), .out(\net10391<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1106.Ivi6  ( .en(GND), .in(\ILAB0102.net25133 ), .out(\ILAB0102.net25699 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0912.Iho1  ( .en(GND), .in(\ILAB0102.net18517 ), .out(\ILAB0102.net18922 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1301.Iho1  ( .en(GND), .in(\net10391<0> ), .out(\ILAB0103.net20452 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0805.Iho1  ( .en(GND), .in(\ILAB0102.net25114 ), .out(\ILAB0102.net17347 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0806.Ivi7  ( .en(GND), .in(\ILAB0102.net25699 ), .out(\ILAB0102.net18634 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0915.Iho2  ( .en(GND), .in(\ILAB0102.net18922 ), .out(\net10407<2> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0608.Ivi7  ( .en(GND), .in(\ILAB0102.net25159 ), .out(\ILAB0102.net19624 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1112.Ivi6  ( .en(GND), .in(\ILAB0102.net16222 ), .out(\ILAB0102.net21379 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1116.Iho2  ( .en(GND), .in(\net10399<0> ), .out(\net10399<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0812.Ivi7  ( .en(GND), .in(\ILAB0102.net21379 ), .out(\ILAB0102.net18679 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0715.Ivi6  ( .en(GND), .in(\ILAB0102.net18922 ), .out(\ILAB0102.net22099 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0903.Ivi7  ( .en(GND), .in(\ILAB0103.net20452 ), .out(\ILAB0103.net20299 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0601.Ivi7  ( .en(GND), .in(\net10407<2> ), .out(\ILAB0103.net20614 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0711.Iho2  ( .en(GND), .in(\ILAB0102.net25159 ), .out(\ILAB0102.net21488 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0814.Iho2  ( .en(GND), .in(\ILAB0102.net16222 ), .out(\ILAB0102.net18878 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0501.Ivo2  ( .en(GND), .in(\ILAB0103.net20614 ), .out(\ILAB0103.net20522 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0905.Iho3  ( .en(GND), .in(\ILAB0102.ILE0905.net2656 ), .out(\ILAB0102.net25404 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0806.Ivo3  ( .en(GND), .in(\ILAB0102.ILE0806.net2656 ), .out(\ILAB0102.net24660 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0710.Iho1  ( .en(GND), .in(\ILAB0102.net24660 ), .out(\ILAB0102.net24142 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0906.Iho1  ( .en(GND), .in(\ILAB0102.net24660 ), .out(\ILAB0102.net24637 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0910.Iho1  ( .en(GND), .in(\ILAB0102.net24637 ), .out(\ILAB0102.net23692 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0906.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0906.net2656 ), .out(\ILAB0102.net24664 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0913.Iho3  ( .en(GND), .in(\ILAB0102.ILE0913.net2656 ), .out(\ILAB0102.net25494 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1014.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1014.net2656 ), .out(\ILAB0102.net23494 ));
  inv_8_UCCLAB \ILAB0102.ILE1014.I666  ( .a(\ILAB0102.ILE1014.net0541 ), .x(\ILAB0102.net21416 ));
  inv_4_UCCLAB \ILAB0102.ILE1115.I714  ( .a(\ILAB0102.net21416 ), .x(\ILAB0102.ILE1115.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0914.Ivo1  ( .en(GND), .in(\ILAB0102.ILE0914.net2656 ), .out(\ILAB0102.net23269 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1115.Iho3  ( .en(GND), .in(\ILAB0102.ILE1115.net2656 ), .out(\ILAB0102.net24504 ));
  inv_8_UCCLAB \ILAB0103.ILE1002.I666  ( .a(\ILAB0103.ILE1002.net0541 ), .x(\ILAB0103.net16556 ));
  inv_4_UCCLAB \ILAB0103.ILE1101.I714  ( .a(\ILAB0103.net16556 ), .x(\ILAB0103.ILE1101.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1116.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1116.net2656 ), .out(\ILAB0102.net21739 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1016.Ivo2  ( .en(GND), .in(\ILAB0102.net21739 ), .out(\ILAB0102.net21197 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1101.Ivo1  ( .en(GND), .in(\ILAB0103.ILE1101.net2656 ), .out(\ILAB0103.net20884 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1202.Ihi7  ( .en(GND), .in(\ILAB0103.ILE1202.net2656 ), .out(\net10395<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1202.Ivi6  ( .en(GND), .in(\ILAB0103.ILE1202.net2656 ), .out(\ILAB0103.net26554 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0902.Ivi7  ( .en(GND), .in(\ILAB0103.net26554 ), .out(\ILAB0103.net26194 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1201.Iho3  ( .en(GND), .in(\ILAB0103.ILE1201.net2656 ), .out(\ILAB0103.net15504 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0901.Ivi7  ( .en(GND), .in(\ILAB0103.ILE0901.net2656 ), .out(\ILAB0103.net20929 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0802.Ihi7  ( .en(GND), .in(\ILAB0103.ILE0802.net2656 ), .out(\net10411<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0802.Ivi7  ( .en(GND), .in(\ILAB0103.ILE0802.net2656 ), .out(\ILAB0103.net26149 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0801.Iho2  ( .en(GND), .in(\net10411<1> ), .out(\ILAB0103.net20678 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0801.Iho3  ( .en(GND), .in(\ILAB0103.ILE0801.net2656 ), .out(\ILAB0103.net20679 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1001.Ihi5  ( .en(GND), .in(\ILAB0103.ILE1001.net2656 ), .out(\net10403<2> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1015.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1015.net2656 ), .out(\ILAB0102.net24484 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1015.Iho3  ( .en(GND), .in(\ILAB0102.ILE1015.net2656 ), .out(\ILAB0102.net24459 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1015.Ivi5  ( .en(GND), .in(\ILAB0102.ILE1015.net2656 ), .out(\ILAB0102.net24482 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0915.Ivo2  ( .en(GND), .in(\ILAB0102.net24484 ), .out(\ILAB0102.net24527 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1016.Ihi7  ( .en(GND), .in(\ILAB0102.ILE1016.net2656 ), .out(\ILAB0102.net21667 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0915.Iho3  ( .en(GND), .in(\ILAB0102.ILE0915.net2656 ), .out(\ILAB0102.net22164 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0902.Ivi5  ( .en(GND), .in(\ILAB0103.ILE0902.net2656 ), .out(\ILAB0103.net26192 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0902.Ihi7  ( .en(GND), .in(\ILAB0103.ILE0902.net2656 ), .out(\net10407<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0916.Iho1  ( .en(GND), .in(\ILAB0102.ILE0916.net2656 ), .out(\net10407<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0816.Ihi7  ( .en(GND), .in(\ILAB0102.ILE0816.net2656 ), .out(\ILAB0102.net18652 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0715.Ivo1  ( .en(GND), .in(\ILAB0102.ILE0715.net2656 ), .out(\ILAB0102.net24529 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0715.Ivi5  ( .en(GND), .in(\ILAB0102.ILE0715.net2656 ), .out(\ILAB0102.net24212 ));
  inv_8_UCCLAB \ILAB0102.ILE0715.I666  ( .a(\ILAB0102.ILE0715.net0541 ), .x(\ILAB0102.net22406 ));
  inv_4_UCCLAB \ILAB0102.ILE0814.I714  ( .a(\ILAB0102.net22406 ), .x(\ILAB0102.ILE0814.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0815.Ivi5  ( .en(GND), .in(\ILAB0102.ILE0815.net2656 ), .out(\ILAB0102.net22097 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0814.Ihi7  ( .en(GND), .in(\ILAB0102.ILE0814.net2656 ), .out(\ILAB0102.net23602 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0810.Ihi5  ( .en(GND), .in(\ILAB0102.ILE0810.net2656 ), .out(\ILAB0102.net17978 ));
  inv_8_UCCLAB \ILAB0102.ILE0810.I666  ( .a(\ILAB0102.ILE0810.net0541 ), .x(\ILAB0102.net17636 ));
  inv_4_UCCLAB \ILAB0102.ILE0711.I712  ( .a(\ILAB0102.net17636 ), .x(\ILAB0102.ILE0711.net0562 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0811.Ihi5  ( .en(GND), .in(\ILAB0102.ILE0811.net2656 ), .out(\ILAB0102.net17618 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0809.Ihi5  ( .en(GND), .in(\ILAB0102.ILE0809.net2656 ), .out(\ILAB0102.net25223 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1007.Ihi6  ( .en(GND), .in(\ILAB0102.ILE1007.net2656 ), .out(\ILAB0102.net23107 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1007.Ivi5  ( .en(GND), .in(\ILAB0102.ILE1007.net2656 ), .out(\ILAB0102.net25832 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0804.Ivi7  ( .en(GND), .in(\ILAB0102.net23107 ), .out(\ILAB0102.net25609 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0907.Ivo3  ( .en(GND), .in(\ILAB0102.ILE0907.net2656 ), .out(\ILAB0102.net25830 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1104.Ihi7  ( .en(GND), .in(\ILAB0102.ILE1104.net2656 ), .out(\net17194<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1102.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1102.net2656 ), .out(\ILAB0102.net26689 ));
  inv_8_UCCLAB \ILAB0102.ILE1102.I666  ( .a(\ILAB0102.ILE1102.net0541 ), .x(\ILAB0102.net16601 ));
  inv_4_UCCLAB \ILAB0102.ILE1003.I712  ( .a(\ILAB0102.net16601 ), .x(\ILAB0102.ILE1003.net0562 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1102.Iho1  ( .en(GND), .in(\ILAB0102.ILE1102.net2656 ), .out(\ILAB0102.net26662 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1103.Ihi7  ( .en(GND), .in(\ILAB0102.ILE1103.net2656 ), .out(\net17194<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1003.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1003.net2656 ), .out(\ILAB0102.net17419 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0902.Iho2  ( .en(GND), .in(\ILAB0102.ILE0902.net2656 ), .out(\ILAB0102.net26168 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0902.Ivi5  ( .en(GND), .in(\ILAB0102.ILE0902.net2656 ), .out(\ILAB0102.net26192 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0702.Ivi6  ( .en(GND), .in(\ILAB0102.net26192 ), .out(\ILAB0102.net26149 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0903.Ihi7  ( .en(GND), .in(\ILAB0102.ILE0903.net2656 ), .out(\net17202<3> ));
  inv_8_UCCLAB \ILAB0102.ILE0904.I666  ( .a(\ILAB0102.ILE0904.net0541 ), .x(\ILAB0102.net20291 ));
  inv_4_UCCLAB \ILAB0102.ILE0803.I710  ( .a(\ILAB0102.net20291 ), .x(\ILAB0102.ILE0803.net0558 ));
  inv_8_UCCLAB \ILAB0102.ILE0703.I666  ( .a(\ILAB0102.ILE0703.net0541 ), .x(\ILAB0102.net26456 ));
  inv_4_UCCLAB \ILAB0102.ILE0604.I712  ( .a(\ILAB0102.net26456 ), .x(\ILAB0102.ILE0604.net0562 ));
  inv_4_UCCLAB \ILAB0102.ILE0804.I714  ( .a(\ILAB0102.net26456 ), .x(\ILAB0102.ILE0804.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0703.Ivo3  ( .en(GND), .in(\ILAB0102.ILE0703.net2656 ), .out(\ILAB0102.net20340 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0803.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0803.net2656 ), .out(\ILAB0102.net20344 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0804.Iho3  ( .en(GND), .in(\ILAB0102.ILE0804.net2656 ), .out(\ILAB0102.net25584 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0705.Iho1  ( .en(GND), .in(\ILAB0102.ILE0705.net2656 ), .out(\ILAB0102.net15817 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0705.Ivo1  ( .en(GND), .in(\ILAB0102.ILE0705.net2656 ), .out(\ILAB0102.net17959 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0705.Iho2  ( .en(GND), .in(\ILAB0102.ILE0705.net2656 ), .out(\ILAB0102.net15818 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0707.Iho3  ( .en(GND), .in(\ILAB0102.net15818 ), .out(\ILAB0102.net17214 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0805.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0805.net2656 ), .out(\ILAB0102.net17374 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0807.Iho3  ( .en(GND), .in(\ILAB0102.ILE0807.net2656 ), .out(\ILAB0102.net25224 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0708.Ivo1  ( .en(GND), .in(\ILAB0102.ILE0708.net2656 ), .out(\ILAB0102.net24799 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0708.Ivi5  ( .en(GND), .in(\ILAB0102.ILE0708.net2656 ), .out(\ILAB0102.net21062 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0808.Ivi5  ( .en(GND), .in(\ILAB0102.ILE0808.net2656 ), .out(\ILAB0102.net18002 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0908.Iho3  ( .en(GND), .in(\ILAB0102.ILE0908.net2656 ), .out(\ILAB0102.net18519 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0910.Ihi6  ( .en(GND), .in(\ILAB0102.ILE0910.net2656 ), .out(\ILAB0102.net25942 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0910.Ivi6  ( .en(GND), .in(\ILAB0102.ILE0910.net2656 ), .out(\ILAB0102.net24889 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0910.Ivo3  ( .en(GND), .in(\ILAB0102.ILE0910.net2656 ), .out(\ILAB0102.net24885 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0909.Iho3  ( .en(GND), .in(\ILAB0102.ILE0909.net2656 ), .out(\ILAB0102.net25314 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1010.Ivo3  ( .en(GND), .in(\ILAB0102.ILE1010.net2656 ), .out(\ILAB0102.net24975 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1210.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1210.net2656 ), .out(\ILAB0102.net24754 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1210.Ivi5  ( .en(GND), .in(\ILAB0102.ILE1210.net2656 ), .out(\ILAB0102.net24752 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1210.Ihi6  ( .en(GND), .in(\ILAB0102.ILE1210.net2656 ), .out(\ILAB0102.net17032 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1110.Ivo1  ( .en(GND), .in(\ILAB0102.ILE1110.net2656 ), .out(\ILAB0102.net24079 ));
  sw_b_v2_inv_UCCLAB \ILAB0202.ILE0105.Iho1  ( .en(GND), .in(\ILAB0202.ILE0105.net2656 ), .out(\ILAB0202.net19732 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1504.Iho1  ( .en(GND), .in(\ILAB0102.ILE1504.net2656 ), .out(\ILAB0102.net16177 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1507.Ihi5  ( .en(GND), .in(\ILAB0102.ILE1507.net2656 ), .out(\ILAB0102.net15728 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1406.Ivo1  ( .en(GND), .in(\ILAB0102.ILE1406.net2656 ), .out(\net18572<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1406.Ivi5  ( .en(GND), .in(\ILAB0102.ILE1406.net2656 ), .out(\ILAB0102.net21152 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1406.Ihi5  ( .en(GND), .in(\ILAB0102.ILE1406.net2656 ), .out(\ILAB0102.net25628 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1506.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1506.net2656 ), .out(\ILAB0102.net18184 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1605.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1605.net2656 ), .out(\ILAB0102.net15889 ));
  inv_8_UCCLAB \ILAB0102.ILE1604.I666  ( .a(\ILAB0102.ILE1604.net0541 ), .x(\ILAB0102.net15476 ));
  buftd4_UCCLAB \ILAB0102.I224  ( .a(\ILAB0102.net15476 ), .en(VDD), .x(\ILAB0102.net27188 ));
  mux2p_2_UCCLAB \ILAB0102.I5605.I0  ( .d0(\ILAB0102.net27188 ), .d1(GND), .s0(GND), .x(\ILAB0102.I5605.net29 ));
  invd16_seth_UCCLAB \ILAB0102.I5605.I1  ( .a(\ILAB0102.I5605.net29 ), .c(VDD), .x(\ILAB0102.Clk_int<3> ));
  mux2d1i_1_P_UCCLAB \ILAB0102.I5366.I81  ( .d0(\ILAB0102.Clk_int<3> ), .d1i(GND), .sl0(GND), .x(\ILAB0102.I5366.net0102 ));
  invd52_UCCLAB \ILAB0102.I5366.I77  ( .a(\ILAB0102.I5366.net0102 ), .x(\ILAB0102.net15299<0> ));
  invd32_UCCLAB \ILAB0102.I5591.I0  ( .a(\ILAB0102.net15299<0> ), .x(\ILAB0102.Clk_LAB<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1505.Ihi6  ( .en(GND), .in(\ILAB0102.ILE1505.net2656 ), .out(\ILAB0102.net26347 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1506.Iho1  ( .en(GND), .in(\ILAB0102.net26347 ), .out(\ILAB0102.net18157 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1506.Ivi5  ( .en(GND), .in(\ILAB0102.net18157 ), .out(\ILAB0102.net18182 ));
  inv_8_UCCLAB \ILAB0102.ILE1406.I666  ( .a(\ILAB0102.net18182 ), .x(\ILAB0102.net25061 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1408.Ivo1  ( .en(GND), .in(\ILAB0102.ILE1408.net2656 ), .out(\net18564<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1408.Ihi5  ( .en(GND), .in(\ILAB0102.ILE1408.net2656 ), .out(\ILAB0102.net21128 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1407.Iho3  ( .en(GND), .in(\ILAB0102.ILE1407.net2656 ), .out(\ILAB0102.net25764 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1508.Iho1  ( .en(GND), .in(\ILAB0102.ILE1508.net2656 ), .out(\ILAB0102.net19552 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1512.Iho1  ( .en(GND), .in(\ILAB0102.net19552 ), .out(\ILAB0102.net19642 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1416.Ivo1  ( .en(GND), .in(\ILAB0102.ILE1416.net2656 ), .out(\net18532<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1416.Ivi5  ( .en(GND), .in(\ILAB0102.ILE1416.net2656 ), .out(\ILAB0102.net17912 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1202.Iho3  ( .en(GND), .in(\ILAB0102.net17912 ), .out(\ILAB0103.net26574 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1516.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1516.net2656 ), .out(\ILAB0102.net18814 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1316.Iho3  ( .en(GND), .in(\ILAB0102.ILE1316.net2656 ), .out(\net10391<4> ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1302.Ihi5  ( .en(GND), .in(\ILAB0103.ILE1302.net2656 ), .out(\net10391<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1302.Ihi7  ( .en(GND), .in(\ILAB0103.ILE1302.net2656 ), .out(\net10391<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1302.Ivi6  ( .en(GND), .in(\ILAB0103.ILE1302.net2656 ), .out(\ILAB0103.net26329 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1301.Iho3  ( .en(GND), .in(\ILAB0103.ILE1301.net2656 ), .out(\ILAB0103.net20454 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1315.Ivo1  ( .en(GND), .in(\ILAB0102.ILE1315.net2656 ), .out(\net18536<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1414.Ivi5  ( .en(GND), .in(\ILAB0102.ILE1414.net2656 ), .out(\ILAB0102.net19847 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1414.Iho1  ( .en(GND), .in(\ILAB0102.ILE1414.net2656 ), .out(\net10387<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1414.Ihi5  ( .en(GND), .in(\ILAB0102.ILE1414.net2656 ), .out(\ILAB0102.net19373 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1412.Ihi6  ( .en(GND), .in(\ILAB0102.net19373 ), .out(\ILAB0102.net18067 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1409.Ihi7  ( .en(GND), .in(\ILAB0102.net18067 ), .out(\ILAB0102.net25042 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1405.Ihi7  ( .en(GND), .in(\ILAB0102.net25042 ), .out(\ILAB0102.net20812 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1405.Ivi7  ( .en(GND), .in(\ILAB0102.net25042 ), .out(\ILAB0102.net25069 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1415.Ihi7  ( .en(GND), .in(\ILAB0102.ILE1415.net2656 ), .out(\ILAB0102.net20407 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1305.Ivo3  ( .en(GND), .in(\ILAB0102.ILE1305.net2656 ), .out(\ILAB0102.net25065 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1404.Iho3  ( .en(GND), .in(\ILAB0102.ILE1404.net2656 ), .out(\ILAB0102.net25629 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1405.Ivi5  ( .en(GND), .in(\ILAB0102.ILE1405.net2656 ), .out(\ILAB0102.net25067 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1205.Ivi6  ( .en(GND), .in(\ILAB0102.net25067 ), .out(\ILAB0102.net15934 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1004.Iho3  ( .en(GND), .in(\ILAB0102.ILE1004.net2656 ), .out(\ILAB0102.net23109 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1004.Ivi5  ( .en(GND), .in(\ILAB0102.ILE1004.net2656 ), .out(\ILAB0102.net23132 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0808.Iho1  ( .en(GND), .in(\ILAB0102.net23132 ), .out(\ILAB0102.net17977 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1004.Ihi7  ( .en(GND), .in(\ILAB0102.ILE1004.net2656 ), .out(\net17198<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1005.Ihi7  ( .en(GND), .in(\ILAB0102.ILE1005.net2656 ), .out(\ILAB0102.net16537 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE1014.Ihi6  ( .en(GND), .in(\ILAB0401.ILE1014.net2656 ), .out(\ILAB0401.net22657 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE1014.Ivi7  ( .en(GND), .in(\ILAB0401.ILE1014.net2656 ), .out(\ILAB0401.net23494 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE1011.Ivi6  ( .en(GND), .in(\ILAB0401.net22657 ), .out(\ILAB0401.net23044 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0710.Ivo1  ( .en(GND), .in(\ILAB0401.ILE0710.net2656 ), .out(\ILAB0401.net24979 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0710.Ivo2  ( .en(GND), .in(\ILAB0401.ILE0710.net2656 ), .out(\ILAB0401.net23717 ));
  inv_8_UCCLAB \ILAB0401.ILE0710.I666  ( .a(\ILAB0401.ILE0710.net0541 ), .x(\ILAB0401.net15656 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0910.Ivo3  ( .en(GND), .in(\ILAB0401.net23717 ), .out(\ILAB0401.net24885 ));
  inv_4_UCCLAB \ILAB0401.ILE0811.I714  ( .a(\ILAB0401.net15656 ), .x(\ILAB0401.ILE0811.net01345 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0710.Iho2  ( .en(GND), .in(\ILAB0401.ILE0710.net2656 ), .out(\ILAB0401.net24143 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0712.Iho3  ( .en(GND), .in(\ILAB0401.net24143 ), .out(\ILAB0401.net19914 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE1010.Ivo2  ( .en(GND), .in(\ILAB0401.net24979 ), .out(\ILAB0401.net24752 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE1012.Iho3  ( .en(GND), .in(\ILAB0401.net24752 ), .out(\ILAB0401.net21669 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0811.Ivi7  ( .en(GND), .in(\ILAB0401.ILE0811.net2656 ), .out(\ILAB0401.net18499 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0711.Ivo2  ( .en(GND), .in(\ILAB0401.net18499 ), .out(\ILAB0401.net18992 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0812.Ivi6  ( .en(GND), .in(\ILAB0401.ILE0812.net2656 ), .out(\ILAB0401.net18949 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0812.Ivi5  ( .en(GND), .in(\ILAB0401.ILE0812.net2656 ), .out(\ILAB0401.net18677 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0613.Iho1  ( .en(GND), .in(\ILAB0401.net18949 ), .out(\net16308<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0512.Ihi6  ( .en(GND), .in(\ILAB0401.net18949 ), .out(\ILAB0401.net19102 ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0601.Iho1  ( .en(GND), .in(\net16308<0> ), .out(\ILAB0402.net20587 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0513.Iho1  ( .en(GND), .in(\ILAB0401.net19102 ), .out(\net16312<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0201.Ivi7  ( .en(GND), .in(\net16312<0> ), .out(\net11344<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE1012.Ivi7  ( .en(GND), .in(\ILAB0401.ILE1012.net2656 ), .out(\ILAB0401.net21694 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0814.Ihi5  ( .en(GND), .in(\ILAB0401.ILE0814.net2656 ), .out(\ILAB0401.net18653 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0814.Ihi6  ( .en(GND), .in(\ILAB0401.ILE0814.net2656 ), .out(\ILAB0401.net18472 ));
  inv_8_UCCLAB \ILAB0401.ILE0814.I666  ( .a(\ILAB0401.ILE0814.net0541 ), .x(\ILAB0401.net22541 ));
  inv_4_UCCLAB \ILAB0401.ILE0713.I711  ( .a(\ILAB0401.net22541 ), .x(\ILAB0401.ILE0713.net0560 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0814.Ivi6  ( .en(GND), .in(\ILAB0401.ILE0814.net2656 ), .out(\ILAB0401.net19174 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0712.Iho2  ( .en(GND), .in(\ILAB0401.ILE0712.net2656 ), .out(\ILAB0401.net19913 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0712.Ihi6  ( .en(GND), .in(\ILAB0401.ILE0712.net2656 ), .out(\ILAB0401.net15637 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0713.Iho1  ( .en(GND), .in(\ILAB0401.net15637 ), .out(\net16304<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0401.Ivi7  ( .en(GND), .in(\net16304<0> ), .out(\net11344<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0302.ILE1601.Ivi7  ( .en(GND), .in(\net11344<6> ), .out(\ILAB0302.net20569 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0415.Ivi7  ( .en(GND), .in(\net16304<0> ), .out(\net16271<6> ));
  inv_8_UCCLAB \ILAB0401.ILE0716.I666  ( .a(\net16304<0> ), .x(\net16244<1> ));
  buf4_12_UCCLAB \ILAB0401.I4397  ( .a(\net16244<1> ), .x(\ILAB0401.net27305 ));
  buftid52C_UCCLAB \ILAB0401.I4462  ( .a(\ILAB0401.net27305 ), .ne(GND), .x(\net8320<7> ));
  inv_4_UCCLAB \ILAB0401.ILE0116.I715  ( .a(\net8320<7> ), .x(\ILAB0401.ILE0116.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0414.Ivo1  ( .en(GND), .in(\ILAB0401.ILE0414.net2656 ), .out(\ILAB0401.net18904 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0516.Ihi7  ( .en(GND), .in(\ILAB0401.ILE0516.net2656 ), .out(\ILAB0401.net19057 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0514.Iho1  ( .en(GND), .in(\ILAB0401.ILE0514.net2656 ), .out(\net16312<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0514.Ivi5  ( .en(GND), .in(\ILAB0401.ILE0514.net2656 ), .out(\ILAB0401.net19802 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0314.Ivi6  ( .en(GND), .in(\ILAB0401.net19802 ), .out(\net16275<6> ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0514.Ivo2  ( .en(GND), .in(\ILAB0401.ILE0514.net2656 ), .out(\ILAB0401.net22412 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0514.Ivi7  ( .en(GND), .in(\ILAB0401.ILE0514.net2656 ), .out(\ILAB0401.net19804 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0515.Ivo1  ( .en(GND), .in(\ILAB0401.ILE0515.net2656 ), .out(\ILAB0401.net22189 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0515.Ihi5  ( .en(GND), .in(\ILAB0401.ILE0515.net2656 ), .out(\ILAB0401.net18293 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0513.Ihi6  ( .en(GND), .in(\ILAB0401.net18293 ), .out(\ILAB0401.net23917 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0115.Ihi7  ( .en(GND), .in(\ILAB0401.ILE0115.net2656 ), .out(\ILAB0401.net23197 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0116.Ivo1  ( .en(GND), .in(\ILAB0401.ILE0116.net2656 ), .out(\ILAB0401.net17014 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0116.Ihi7  ( .en(GND), .in(\ILAB0401.ILE0116.net2656 ), .out(\ILAB0401.net21892 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0116.Ihi5  ( .en(GND), .in(\ILAB0401.ILE0116.net2656 ), .out(\ILAB0401.net23648 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0114.Ihi7  ( .en(GND), .in(\ILAB0401.ILE0114.net2656 ), .out(\ILAB0401.net25267 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0412.Ivo1  ( .en(GND), .in(\ILAB0401.ILE0412.net2656 ), .out(\ILAB0401.net18679 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0513.Ihi5  ( .en(GND), .in(\ILAB0401.ILE0513.net2656 ), .out(\ILAB0401.net20363 ));
  inv_8_UCCLAB \ILAB0401.ILE0513.I666  ( .a(\ILAB0401.ILE0513.net0541 ), .x(\ILAB0401.net19076 ));
  inv_4_UCCLAB \ILAB0401.ILE0612.I713  ( .a(\ILAB0401.net19076 ), .x(\ILAB0401.ILE0612.net01342 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0513.Ivo3  ( .en(GND), .in(\ILAB0401.ILE0513.net2656 ), .out(\ILAB0401.net19350 ));
  inv_8_UCCLAB \ILAB0401.ILE0613.I666  ( .a(\ILAB0401.ILE0613.net0541 ), .x(\ILAB0401.net19706 ));
  inv_4_UCCLAB \ILAB0401.ILE0714.I715  ( .a(\ILAB0401.net19706 ), .x(\ILAB0401.ILE0714.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0613.Iho2  ( .en(GND), .in(\ILAB0401.ILE0613.net2656 ), .out(\ILAB0401.net19328 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0615.Iho3  ( .en(GND), .in(\ILAB0401.net19328 ), .out(\ILAB0401.net23964 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0612.Ivi7  ( .en(GND), .in(\ILAB0401.ILE0612.net2656 ), .out(\ILAB0401.net19714 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0512.Ivi7  ( .en(GND), .in(\ILAB0401.ILE0512.net2656 ), .out(\ILAB0401.net19084 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0212.Ivo3  ( .en(GND), .in(\ILAB0401.ILE0212.net2656 ), .out(\ILAB0401.net24930 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0214.Ihi7  ( .en(GND), .in(\ILAB0401.ILE0214.net2656 ), .out(\ILAB0401.net25537 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0213.Ivo3  ( .en(GND), .in(\ILAB0401.ILE0213.net2656 ), .out(\ILAB0401.net23175 ));
  inv_8_UCCLAB \ILAB0402.ILE0701.I666  ( .a(\ILAB0402.ILE0701.net0541 ), .x(\net16244<0> ));
  inv_4_UCCLAB \ILAB0401.ILE0616.I710  ( .a(\net16244<0> ), .x(\ILAB0401.ILE0616.net0558 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0315.Iho1  ( .en(GND), .in(\ILAB0401.ILE0315.net2656 ), .out(\net16320<3> ));
  inv_8_UCCLAB \ILAB0401.ILE0315.I666  ( .a(\ILAB0401.ILE0315.net0541 ), .x(\ILAB0401.net23801 ));
  inv_4_UCCLAB \ILAB0401.ILE0416.I713  ( .a(\ILAB0401.net23801 ), .x(\ILAB0401.ILE0416.net01342 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0315.Ivo3  ( .en(GND), .in(\ILAB0401.ILE0315.net2656 ), .out(\ILAB0401.net22365 ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0301.Ihi5  ( .en(GND), .in(\ILAB0402.ILE0301.net2656 ), .out(\net16320<2> ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0415.Ihi5  ( .en(GND), .in(\ILAB0401.ILE0415.net2656 ), .out(\ILAB0401.net26078 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0415.Ihi7  ( .en(GND), .in(\ILAB0401.ILE0415.net2656 ), .out(\ILAB0401.net19867 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0414.Iho2  ( .en(GND), .in(\ILAB0401.net19867 ), .out(\ILAB0401.net19238 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0614.Iho3  ( .en(GND), .in(\ILAB0401.ILE0614.net2656 ), .out(\ILAB0401.net22119 ));
  inv_8_UCCLAB \ILAB0401.ILE0614.I666  ( .a(\ILAB0401.ILE0614.net0541 ), .x(\ILAB0401.net19346 ));
  inv_4_UCCLAB \ILAB0401.ILE0715.I715  ( .a(\ILAB0401.net19346 ), .x(\ILAB0401.ILE0715.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0715.Ihi7  ( .en(GND), .in(\ILAB0401.ILE0715.net2656 ), .out(\ILAB0401.net21487 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0714.Iho2  ( .en(GND), .in(\ILAB0401.net21487 ), .out(\ILAB0401.net22388 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0715.Iho1  ( .en(GND), .in(\ILAB0401.ILE0715.net2656 ), .out(\net16304<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0302.Ivi7  ( .en(GND), .in(\net16304<3> ), .out(\net11340<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0615.Iho1  ( .en(GND), .in(\ILAB0401.ILE0615.net2656 ), .out(\net16308<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0615.Iho2  ( .en(GND), .in(\ILAB0401.ILE0615.net2656 ), .out(\net16308<2> ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0316.Ivi7  ( .en(GND), .in(\ILAB0401.ILE0316.net2656 ), .out(\net16267<3> ));
  inv_8_UCCLAB \ILAB0401.ILE0316.I666  ( .a(\ILAB0401.ILE0316.net0541 ), .x(\net16248<1> ));
  inv_4_UCCLAB \ILAB0402.ILE0401.I713  ( .a(\net16248<1> ), .x(\ILAB0402.ILE0401.net01342 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0416.Ivo1  ( .en(GND), .in(\ILAB0401.ILE0416.net2656 ), .out(\ILAB0401.net17464 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0616.Ivo1  ( .en(GND), .in(\ILAB0401.ILE0616.net2656 ), .out(\ILAB0401.net21604 ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0501.Ivo1  ( .en(GND), .in(\ILAB0402.ILE0501.net2656 ), .out(\ILAB0402.net20929 ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0401.Ivo2  ( .en(GND), .in(\ILAB0402.ILE0401.net2656 ), .out(\ILAB0402.net20612 ));
  inv_8_UCCLAB \ILAB0402.ILE0601.I666  ( .a(\ILAB0402.ILE0601.net0541 ), .x(\net16245<0> ));
  inv_4_UCCLAB \ILAB0402.ILE0502.I712  ( .a(\net16245<0> ), .x(\ILAB0402.ILE0502.net0562 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0216.Iho3  ( .en(GND), .in(\ILAB0401.ILE0216.net2656 ), .out(\net16324<4> ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0201.Iho3  ( .en(GND), .in(\ILAB0402.ILE0201.net2656 ), .out(\ILAB0402.net16944 ));
  sw_b_v2_inv_UCCLAB \ILAB0402.ILE0101.Iho3  ( .en(GND), .in(\ILAB0402.ILE0101.net2656 ), .out(\ILAB0402.net16719 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1302.Ivi5  ( .en(GND), .in(\ILAB0102.ILE1302.net2656 ), .out(\ILAB0102.net26552 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1102.Ivi6  ( .en(GND), .in(\ILAB0102.net26552 ), .out(\ILAB0102.net26599 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0901.Ihi7  ( .en(GND), .in(\ILAB0102.ILE0901.net2656 ), .out(\net17202<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0911.Ihi5  ( .en(GND), .in(\ILAB0401.ILE0911.net2656 ), .out(\ILAB0401.net25313 ));
  inv_8_UCCLAB \ILAB0401.ILE0911.I666  ( .a(\ILAB0401.ILE0911.net0541 ), .x(\ILAB0401.net23711 ));
  inv_4_UCCLAB \ILAB0401.ILE1010.I713  ( .a(\ILAB0401.net23711 ), .x(\ILAB0401.ILE1010.net01342 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0911.Ivo3  ( .en(GND), .in(\ILAB0401.ILE0911.net2656 ), .out(\ILAB0401.net22680 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0911.Iho2  ( .en(GND), .in(\ILAB0401.ILE0911.net2656 ), .out(\ILAB0401.net18968 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0913.Iho3  ( .en(GND), .in(\ILAB0401.net18968 ), .out(\ILAB0401.net25494 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE1013.Ivi7  ( .en(GND), .in(\ILAB0401.ILE1013.net2656 ), .out(\ILAB0401.net21424 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0613.Ivi7  ( .en(GND), .in(\ILAB0401.net21424 ), .out(\ILAB0401.net19354 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0213.Ivi7  ( .en(GND), .in(\ILAB0401.net19354 ), .out(\net16279<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0301.ILE1413.Ivi7  ( .en(GND), .in(\net16279<1> ), .out(\ILAB0301.net18364 ));
  sw_b_v2_inv_UCCLAB \ILAB0301.ILE1013.Ivi7  ( .en(GND), .in(\ILAB0301.net18364 ), .out(\ILAB0301.net21424 ));
  sw_b_v2_inv_UCCLAB \ILAB0301.ILE0613.Ivi7  ( .en(GND), .in(\ILAB0301.net21424 ), .out(\ILAB0301.net19354 ));
  sw_b_v2_inv_UCCLAB \ILAB0301.ILE0213.Ivi7  ( .en(GND), .in(\ILAB0301.net19354 ), .out(\net16430<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0201.ILE1413.Ivi7  ( .en(GND), .in(\net16430<1> ), .out(\ILAB0201.net18364 ));
  sw_b_v2_inv_UCCLAB \ILAB0201.ILE1013.Ivi7  ( .en(GND), .in(\ILAB0201.net18364 ), .out(\ILAB0201.net21424 ));
  sw_b_v2_inv_UCCLAB \ILAB0201.ILE0613.Ivi7  ( .en(GND), .in(\ILAB0201.net21424 ), .out(\ILAB0201.net19354 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE1010.Ivi7  ( .en(GND), .in(\ILAB0401.ILE1010.net2656 ), .out(\ILAB0401.net24889 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0910.Ivo2  ( .en(GND), .in(\ILAB0401.net24889 ), .out(\ILAB0401.net24977 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0912.Iho3  ( .en(GND), .in(\ILAB0401.ILE0912.net2656 ), .out(\ILAB0401.net18924 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0912.Iho1  ( .en(GND), .in(\ILAB0401.ILE0912.net2656 ), .out(\ILAB0401.net18922 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0913.Ivi7  ( .en(GND), .in(\ILAB0401.ILE0913.net2656 ), .out(\ILAB0401.net25519 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0713.Ivo1  ( .en(GND), .in(\ILAB0401.ILE0713.net2656 ), .out(\ILAB0401.net21559 ));
  inv_8_UCCLAB \ILAB0401.ILE0714.I666  ( .a(\ILAB0401.ILE0714.net0541 ), .x(\ILAB0401.net19976 ));
  inv_4_UCCLAB \ILAB0401.ILE0813.I715  ( .a(\ILAB0401.net19976 ), .x(\ILAB0401.ILE0813.net01339 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0813.Iho3  ( .en(GND), .in(\ILAB0401.ILE0813.net2656 ), .out(\ILAB0401.net22524 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE1011.Ivi7  ( .en(GND), .in(\ILAB0401.ILE1011.net2656 ), .out(\ILAB0401.net22684 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0911.Ivo2  ( .en(GND), .in(\ILAB0401.net22684 ), .out(\ILAB0401.net23042 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0914.Ivo1  ( .en(GND), .in(\ILAB0401.ILE0914.net2656 ), .out(\ILAB0401.net23269 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0910.Ivi7  ( .en(GND), .in(\ILAB0401.ILE0910.net2656 ), .out(\ILAB0401.net23719 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0611.Ivi6  ( .en(GND), .in(\ILAB0401.ILE0611.net2656 ), .out(\ILAB0401.net21514 ));
  inv_8_UCCLAB \ILAB0401.ILE0810.I666  ( .a(\ILAB0401.ILE0810.net0541 ), .x(\ILAB0401.net17636 ));
  inv_4_UCCLAB \ILAB0401.ILE0711.I710  ( .a(\ILAB0401.net17636 ), .x(\ILAB0401.ILE0711.net0558 ));
  sw_b_v2_inv_UCCLAB \ILAB0401.ILE0711.Ihi7  ( .en(GND), .in(\ILAB0401.ILE0711.net2656 ), .out(\ILAB0401.net17212 ));
  sw_b_v2_inv_UCCLAB \ILAB0201.ILE0313.Iho3  ( .en(GND), .in(\ILAB0201.ILE0313.net2656 ), .out(\ILAB0201.net23154 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0503.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0503.net2656 ), .out(\Fast_out_28<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0713.Iho3  ( .en(GND), .in(\ILAB0102.ILE0713.net2656 ), .out(\ILAB0102.net19959 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0615.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0615.net2656 ), .out(\ILAB0102.net23989 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1003.Iho3  ( .en(GND), .in(\ILAB0103.ILE1003.net2656 ), .out(\ILAB0103.net17394 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0702.Ivi7  ( .en(GND), .in(\ILAB0103.ILE0702.net2656 ), .out(\ILAB0103.net26464 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0502.Iho3  ( .en(GND), .in(\ILAB0103.ILE0502.net2656 ), .out(\ILAB0103.net26259 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0903.Iho3  ( .en(GND), .in(\ILAB0103.ILE0903.net2656 ), .out(\ILAB0103.net20274 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0703.Iho3  ( .en(GND), .in(\ILAB0103.ILE0703.net2656 ), .out(\ILAB0103.net15684 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0501.Ivi7  ( .en(GND), .in(\ILAB0103.ILE0501.net2656 ), .out(\Fast_out_29<7> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0711.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0711.net2656 ), .out(\ILAB0102.net21514 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0504.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0504.net2656 ), .out(\Fast_out_28<4> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0802.Ihi7  ( .en(GND), .in(\ILAB0102.ILE0802.net2656 ), .out(\net17206<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0602.Ihi5  ( .en(GND), .in(\ILAB0102.ILE0602.net2656 ), .out(\net17214<5> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0604.Iho3  ( .en(GND), .in(\ILAB0102.ILE0604.net2656 ), .out(\ILAB0102.net25989 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0706.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0706.net2656 ), .out(\ILAB0102.net16069 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0608.Ivi5  ( .en(GND), .in(\ILAB0102.ILE0608.net2656 ), .out(\ILAB0102.net19622 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0710.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0710.net2656 ), .out(\ILAB0102.net24169 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1011.Iho3  ( .en(GND), .in(\ILAB0102.ILE1011.net2656 ), .out(\ILAB0102.net22659 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1306.Iho3  ( .en(GND), .in(\ILAB0102.ILE1306.net2656 ), .out(\ILAB0102.net18699 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1312.Ivi7  ( .en(GND), .in(\ILAB0102.ILE1312.net2656 ), .out(\ILAB0102.net21244 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1203.Iho3  ( .en(GND), .in(\ILAB0103.ILE1203.net2656 ), .out(\ILAB0103.net15594 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE1102.Iho3  ( .en(GND), .in(\ILAB0103.ILE1102.net2656 ), .out(\ILAB0103.net26664 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE1215.Iho3  ( .en(GND), .in(\ILAB0102.ILE1215.net2656 ), .out(\ILAB0102.net24414 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0812.Iho3  ( .en(GND), .in(\ILAB0102.ILE0812.net2656 ), .out(\ILAB0102.net18654 ));
  sw_b_v2_inv_UCCLAB \ILAB0302.ILE1601.Ivi6  ( .en(GND), .in(\ILAB0302.ILE1601.net2656 ), .out(\net11344<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0308.Ivo1  ( .en(GND), .in(\ILAB0102.ILE0308.net2656 ), .out(\ILAB0102.net21064 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0408.Iho1  ( .en(GND), .in(\ILAB0102.ILE0408.net2656 ), .out(\ILAB0102.net19417 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0716.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0716.net2656 ), .out(\ILAB0102.net19309 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0616.Ihi7  ( .en(GND), .in(\ILAB0102.ILE0616.net2656 ), .out(\ILAB0102.net19687 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0516.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0516.net2656 ), .out(\ILAB0102.net17014 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0416.Ihi5  ( .en(GND), .in(\ILAB0102.ILE0416.net2656 ), .out(\ILAB0102.net19238 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0414.Ihi6  ( .en(GND), .in(\ILAB0102.net19238 ), .out(\ILAB0102.net19867 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0202.Iho3  ( .en(GND), .in(\ILAB0102.ILE0202.net2656 ), .out(\ILAB0102.net26754 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0203.Iho1  ( .en(GND), .in(\ILAB0102.ILE0203.net2656 ), .out(\ILAB0102.net23827 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0207.Iho1  ( .en(GND), .in(\ILAB0102.net23827 ), .out(\ILAB0102.net16852 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0211.Iho1  ( .en(GND), .in(\ILAB0102.net16852 ), .out(\ILAB0102.net23287 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0406.Ivi6  ( .en(GND), .in(\ILAB0102.ILE0406.net2656 ), .out(\Fast_out_28<2> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0506.Iho3  ( .en(GND), .in(\ILAB0102.ILE0506.net2656 ), .out(\ILAB0102.net18744 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0305.Ivo1  ( .en(GND), .in(\ILAB0102.ILE0305.net2656 ), .out(\ILAB0102.net15844 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0405.Iho2  ( .en(GND), .in(\ILAB0102.ILE0405.net2656 ), .out(\ILAB0102.net17753 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0403.Ihi7  ( .en(GND), .in(\ILAB0103.ILE0403.net2656 ), .out(\net10427<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0402.Ihi7  ( .en(GND), .in(\ILAB0103.ILE0402.net2656 ), .out(\net10427<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0414.Ihi7  ( .en(GND), .in(\net10427<1> ), .out(\ILAB0102.net23872 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0604.Iho3  ( .en(GND), .in(\ILAB0103.ILE0604.net2656 ), .out(\ILAB0103.net25989 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0605.Ivi7  ( .en(GND), .in(\ILAB0103.ILE0605.net2656 ), .out(\ILAB0103.net15799 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0401.Iho3  ( .en(GND), .in(\ILAB0102.ILE0401.net2656 ), .out(\ILAB0102.net20724 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0402.Ihi6  ( .en(GND), .in(\ILAB0102.ILE0402.net2656 ), .out(\net17222<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0403.Iho1  ( .en(GND), .in(\net17222<3> ), .out(\ILAB0102.net20182 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0501.Iho3  ( .en(GND), .in(\ILAB0102.ILE0501.net2656 ), .out(\ILAB0102.net20634 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0502.Iho1  ( .en(GND), .in(\ILAB0102.ILE0502.net2656 ), .out(\ILAB0102.net26257 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0505.Iho2  ( .en(GND), .in(\ILAB0102.net26257 ), .out(\ILAB0102.net25448 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0204.Ivo1  ( .en(GND), .in(\ILAB0102.ILE0204.net2656 ), .out(\ILAB0102.net26014 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0304.Iho1  ( .en(GND), .in(\ILAB0102.ILE0304.net2656 ), .out(\ILAB0102.net16132 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0308.Iho1  ( .en(GND), .in(\ILAB0102.net16132 ), .out(\ILAB0102.net15367 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0303.Ihi7  ( .en(GND), .in(\ILAB0103.ILE0303.net2656 ), .out(\net10431<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0302.Ihi7  ( .en(GND), .in(\ILAB0103.ILE0302.net2656 ), .out(\net10431<1> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0514.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0514.net2656 ), .out(\ILAB0102.net19804 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0414.Ihi5  ( .en(GND), .in(\ILAB0102.ILE0414.net2656 ), .out(\ILAB0102.net19013 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0310.Ivo3  ( .en(GND), .in(\ILAB0102.ILE0310.net2656 ), .out(\ILAB0102.net23895 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0410.Iho3  ( .en(GND), .in(\ILAB0102.ILE0410.net2656 ), .out(\ILAB0102.net23874 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0411.Ihi5  ( .en(GND), .in(\ILAB0102.ILE0411.net2656 ), .out(\ILAB0102.net18383 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0409.Ihi6  ( .en(GND), .in(\ILAB0102.net18383 ), .out(\ILAB0102.net18112 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0407.Iho1  ( .en(GND), .in(\ILAB0102.ILE0407.net2656 ), .out(\ILAB0102.net16672 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0404.Ivi6  ( .en(GND), .in(\ILAB0103.ILE0404.net2656 ), .out(\Fast_out_29<4> ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0504.Iho3  ( .en(GND), .in(\ILAB0103.ILE0504.net2656 ), .out(\ILAB0103.net24999 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0804.Iho3  ( .en(GND), .in(\ILAB0103.ILE0804.net2656 ), .out(\ILAB0103.net25584 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0805.Ivi7  ( .en(GND), .in(\ILAB0103.ILE0805.net2656 ), .out(\ILAB0103.net17374 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0612.Ivo3  ( .en(GND), .in(\ILAB0102.ILE0612.net2656 ), .out(\ILAB0102.net19935 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0712.Ihi6  ( .en(GND), .in(\ILAB0102.ILE0712.net2656 ), .out(\ILAB0102.net15637 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0713.Iho1  ( .en(GND), .in(\ILAB0102.net15637 ), .out(\net10415<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0701.Iho1  ( .en(GND), .in(\net10415<0> ), .out(\ILAB0103.net20497 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0705.Ivi7  ( .en(GND), .in(\ILAB0103.ILE0705.net2656 ), .out(\ILAB0103.net15844 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0505.Ihi7  ( .en(GND), .in(\ILAB0103.ILE0505.net2656 ), .out(\ILAB0103.net20632 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0501.Ihi7  ( .en(GND), .in(\ILAB0103.net20632 ), .out(\net10423<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0513.Ihi7  ( .en(GND), .in(\net10423<0> ), .out(\ILAB0102.net19102 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0509.Ihi7  ( .en(GND), .in(\ILAB0102.net19102 ), .out(\ILAB0102.net25447 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0511.Ihi7  ( .en(GND), .in(\ILAB0102.ILE0511.net2656 ), .out(\ILAB0102.net16762 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0510.Ihi5  ( .en(GND), .in(\ILAB0102.ILE0510.net2656 ), .out(\ILAB0102.net19463 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0707.Ivi6  ( .en(GND), .in(\ILAB0102.ILE0707.net2656 ), .out(\ILAB0102.net25249 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0607.Ivi5  ( .en(GND), .in(\ILAB0102.ILE0607.net2656 ), .out(\ILAB0102.net17102 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0507.Iho2  ( .en(GND), .in(\ILAB0102.ILE0507.net2656 ), .out(\ILAB0102.net16763 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0509.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0509.net2656 ), .out(\ILAB0102.net19129 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0409.Ivi5  ( .en(GND), .in(\ILAB0102.ILE0409.net2656 ), .out(\ILAB0102.net18407 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0213.Ivo3  ( .en(GND), .in(\ILAB0102.ILE0213.net2656 ), .out(\ILAB0102.net23175 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0313.Ivo3  ( .en(GND), .in(\ILAB0102.ILE0313.net2656 ), .out(\ILAB0102.net26100 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0413.Ihi5  ( .en(GND), .in(\ILAB0102.ILE0413.net2656 ), .out(\ILAB0102.net19868 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0412.Ivi6  ( .en(GND), .in(\ILAB0102.ILE0412.net2656 ), .out(\ILAB0102.net19084 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0316.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0316.net2656 ), .out(\ELLR15_28<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0216.Ihi7  ( .en(GND), .in(\ILAB0102.ILE0216.net2656 ), .out(\ILAB0102.net22297 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0215.Ivi6  ( .en(GND), .in(\ILAB0102.ILE0215.net2656 ), .out(\ELLR14_28<3> ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0201.Ivo3  ( .en(GND), .in(\ILAB0103.ILE0201.net2656 ), .out(\ILAB0103.net17865 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0301.Ihi7  ( .en(GND), .in(\ILAB0103.ILE0301.net2656 ), .out(\net10431<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0315.Ihi7  ( .en(GND), .in(\ILAB0102.ILE0315.net2656 ), .out(\ILAB0102.net23377 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0513.Ivo1  ( .en(GND), .in(\ILAB0102.ILE0513.net2656 ), .out(\ILAB0102.net25519 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0613.Iho3  ( .en(GND), .in(\ILAB0102.ILE0613.net2656 ), .out(\ILAB0102.net19329 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0701.Ivi7  ( .en(GND), .in(\ILAB0103.ILE0701.net2656 ), .out(\ILAB0103.net20524 ));
  sw_b_v2_inv_UCCLAB \ILAB0103.ILE0601.Ihi7  ( .en(GND), .in(\ILAB0103.ILE0601.net2656 ), .out(\net10419<0> ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0614.Ivi7  ( .en(GND), .in(\ILAB0102.ILE0614.net2656 ), .out(\ILAB0102.net22144 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0311.Iho3  ( .en(GND), .in(\ILAB0102.ILE0311.net2656 ), .out(\ILAB0102.net23379 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0312.Ihi5  ( .en(GND), .in(\ILAB0102.ILE0312.net2656 ), .out(\ILAB0102.net25898 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0310.Ihi6  ( .en(GND), .in(\ILAB0102.net25898 ), .out(\ILAB0102.net25852 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0309.Ihi6  ( .en(GND), .in(\ILAB0102.ILE0309.net2656 ), .out(\ILAB0102.net17527 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0306.Ihi7  ( .en(GND), .in(\ILAB0102.net17527 ), .out(\ILAB0102.net26797 ));
  sw_b_v2_inv_UCCLAB \ILAB0102.ILE0302.Ihi7  ( .en(GND), .in(\ILAB0102.net26797 ), .out(\net17226<1> ));
endmodule
///////////////////////////////////////////////////////
