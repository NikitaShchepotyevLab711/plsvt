module adc7710_wrap (
    input wire clk,
    input wire rst_l,

    // SPI signals //

    inout  wire SDATA,
    input  wire DRDY,
    output wire RFS,
    output wire TFS,
    output wire A0,
    output wire SCLK


);
    
endmodule